module Add(
  input        enable, // @[\\src\\main\\scala\\fpu8\\Add.scala 9:18]
  input  [7:0] a_data, // @[\\src\\main\\scala\\fpu8\\Add.scala 10:13]
  input  [7:0] b_data, // @[\\src\\main\\scala\\fpu8\\Add.scala 11:13]
  input        subtract, // @[\\src\\main\\scala\\fpu8\\Add.scala 12:20]
  input  [1:0] roundingMode, // @[\\src\\main\\scala\\fpu8\\Add.scala 13:24]
  output       sign, // @[\\src\\main\\scala\\fpu8\\Add.scala 14:16]
  output [4:0] exponent, // @[\\src\\main\\scala\\fpu8\\Add.scala 15:20]
  output [3:0] fraction, // @[\\src\\main\\scala\\fpu8\\Add.scala 16:20]
  output       overflow, // @[\\src\\main\\scala\\fpu8\\Add.scala 17:20]
  output       is0, // @[\\src\\main\\scala\\fpu8\\Add.scala 19:15]
  output       isNaN // @[\\src\\main\\scala\\fpu8\\Add.scala 20:17]
);
  wire  compare = a_data[6:0] > b_data[6:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 29:77]
  wire [7:0] greaterOperand_data = compare ? a_data : b_data; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 129:29]
  wire [7:0] smallerOperand_data = compare ? b_data : a_data; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 130:29]
  wire  resultSign = compare ? a_data[7] : b_data[7] ^ subtract; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 131:19]
  wire  subtraction = subtract ^ greaterOperand_data[7] ^ smallerOperand_data[7]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 132:54]
  wire [3:0] exponent_1 = greaterOperand_data[6:3]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 25:28]
  wire  _greaterOperandFraction_T_1 = exponent_1 == 4'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 33:39]
  wire  _greaterOperandFraction_T_2 = ~_greaterOperandFraction_T_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 134:38]
  wire  _smallerOperandFraction_T_1 = smallerOperand_data[6:3] == 4'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 33:39]
  wire  _smallerOperandFraction_T_2 = ~_smallerOperandFraction_T_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 135:38]
  wire  isOnlySmallerDenormalized = _greaterOperandFraction_T_2 & _smallerOperandFraction_T_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 136:60]
  wire [3:0] _shift_T_2 = exponent_1 - 4'h1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 139:31]
  wire [3:0] _shift_T_6 = exponent_1 - smallerOperand_data[6:3]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 140:31]
  wire [3:0] shift = isOnlySmallerDenormalized ? _shift_T_2 : _shift_T_6; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 137:20]
  wire  _shiftedFraction_shifted_T = shift >= 4'h6; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 145:15]
  wire [9:0] _shiftedFraction_shifted_T_1 = {6'h0,_smallerOperandFraction_T_2,smallerOperand_data[2:0]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 146:12]
  wire [9:0] _shiftedFraction_shifted_T_2 = {_smallerOperandFraction_T_2,smallerOperand_data[2:0],6'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 147:12]
  wire [9:0] _shiftedFraction_shifted_T_3 = _shiftedFraction_shifted_T_2 >> shift; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 147:54]
  wire [9:0] shiftedFraction_shifted = _shiftedFraction_shifted_T ? _shiftedFraction_shifted_T_1 :
    _shiftedFraction_shifted_T_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 144:24]
  wire [6:0] smallerOperandFraction_1 = {shiftedFraction_shifted[9:4],|shiftedFraction_shifted[3:0]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 149:10]
  wire [6:0] greaterOperandFraction_1 = {_greaterOperandFraction_T_2,greaterOperand_data[2:0],3'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 151:45]
  wire  _isResultNaN_T_1 = a_data[6:3] == 4'hf; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 35:41]
  wire  _isResultNaN_T_3 = a_data[2:0] == 3'h7; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 39:46]
  wire  _isResultNaN_T_4 = _isResultNaN_T_1 & _isResultNaN_T_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 41:30]
  wire  _isResultNaN_T_6 = b_data[6:3] == 4'hf; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 35:41]
  wire  _isResultNaN_T_8 = b_data[2:0] == 3'h7; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 39:46]
  wire  _isResultNaN_T_9 = _isResultNaN_T_6 & _isResultNaN_T_8; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 41:30]
  wire  isResultNaN = _isResultNaN_T_4 | _isResultNaN_T_9; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 413:37]
  wire  _isResult0_T_2 = a_data[6:0] == b_data[6:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 31:77]
  wire  isResult0 = _isResult0_T_2 & subtraction & ~isResultNaN; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 421:85]
  wire [7:0] _calculatedValue_T_1 = greaterOperandFraction_1 - smallerOperandFraction_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 426:32]
  wire [7:0] _calculatedValue_T_3 = greaterOperandFraction_1 + smallerOperandFraction_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 427:32]
  wire [7:0] calculatedValue = subtraction ? _calculatedValue_T_1 : _calculatedValue_T_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 425:32]
  wire [6:0] _leadingZeros_T_17 = {calculatedValue[0],calculatedValue[1],calculatedValue[2],calculatedValue[3],
    calculatedValue[4],calculatedValue[5],calculatedValue[6]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 58:44]
  wire [2:0] _leadingZeros_T_25 = _leadingZeros_T_17[5] ? 3'h5 : 3'h6; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] _leadingZeros_T_26 = _leadingZeros_T_17[4] ? 3'h4 : _leadingZeros_T_25; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] _leadingZeros_T_27 = _leadingZeros_T_17[3] ? 3'h3 : _leadingZeros_T_26; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] _leadingZeros_T_28 = _leadingZeros_T_17[2] ? 3'h2 : _leadingZeros_T_27; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] _leadingZeros_T_29 = _leadingZeros_T_17[1] ? 3'h1 : _leadingZeros_T_28; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] shift_1 = _leadingZeros_T_17[0] ? 3'h0 : _leadingZeros_T_29; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [7:0] _shiftedValue_T_3 = {calculatedValue[6:0], 1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 63:23]
  wire [8:0] _shiftedValue_T_5 = {calculatedValue[6:0], 2'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 63:23]
  wire [9:0] _shiftedValue_T_7 = {calculatedValue[6:0], 3'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 63:23]
  wire [10:0] _shiftedValue_T_9 = {calculatedValue[6:0], 4'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 63:23]
  wire [11:0] _shiftedValue_T_11 = {calculatedValue[6:0], 5'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 63:23]
  wire [12:0] _shiftedValue_T_13 = {calculatedValue[6:0], 6'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 63:23]
  wire [6:0] _shiftedValue_T_18 = 3'h1 == shift_1 ? _shiftedValue_T_3[6:0] : calculatedValue[6:0]; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [6:0] _shiftedValue_T_20 = 3'h2 == shift_1 ? _shiftedValue_T_5[6:0] : _shiftedValue_T_18; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [6:0] _shiftedValue_T_22 = 3'h3 == shift_1 ? _shiftedValue_T_7[6:0] : _shiftedValue_T_20; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [6:0] _shiftedValue_T_24 = 3'h4 == shift_1 ? _shiftedValue_T_9[6:0] : _shiftedValue_T_22; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [6:0] _shiftedValue_T_26 = 3'h5 == shift_1 ? _shiftedValue_T_11[6:0] : _shiftedValue_T_24; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [6:0] shiftedCalcValue = 3'h6 == shift_1 ? _shiftedValue_T_13[6:0] : _shiftedValue_T_26; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _T_1 = &exponent_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 275:19]
  wire [3:0] _tempExponent_T_1 = exponent_1 + 4'h1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 279:32]
  wire [6:0] _tempFraction_T_3 = {calculatedValue[7:2],|calculatedValue[1:0]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 280:26]
  wire [3:0] _GEN_14 = {{1'd0}, shift_1}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 281:25]
  wire [3:0] _tempExponent_T_3 = exponent_1 - _GEN_14; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 282:32]
  wire [21:0] _GEN_5 = {{15'd0}, calculatedValue[6:0]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 287:47]
  wire [21:0] _tempFraction_T_7 = _GEN_5 << _shift_T_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 287:47]
  wire [21:0] _GEN_0 = exponent_1 > 4'h0 ? _tempFraction_T_7 : {{15'd0}, calculatedValue[6:0]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 286:28 287:22 289:22]
  wire [3:0] _GEN_1 = exponent_1 > _GEN_14 & shiftedCalcValue[6] ? _tempExponent_T_3 : 4'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 281:57 282:20 285:20]
  wire [21:0] _GEN_2 = exponent_1 > _GEN_14 & shiftedCalcValue[6] ? {{15'd0}, shiftedCalcValue} : _GEN_0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 281:57 283:20]
  wire [3:0] _GEN_3 = ~_T_1 & calculatedValue[7] ? _tempExponent_T_1 : _GEN_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 278:54 279:20]
  wire [21:0] _GEN_4 = ~_T_1 & calculatedValue[7] ? {{15'd0}, _tempFraction_T_3} : _GEN_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 278:54 280:20]
  wire [3:0] tempExponent = &exponent_1 & calculatedValue[7] ? exponent_1 : _GEN_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 275:47 276:20]
  wire [21:0] _GEN_6 = &exponent_1 & calculatedValue[7] ? 22'h7f : _GEN_4; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 275:47 277:20]
  wire [6:0] tempFraction = _GEN_6[6:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 273:28]
  wire  _addOne_T_2 = roundingMode == 2'h0 & tempFraction[2]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 234:42]
  wire  _addOne_T_17 = _addOne_T_2 & ~tempFraction[1] & ~tempFraction[0] & tempFraction[3]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 235:90]
  wire  _addOne_T_18 = roundingMode == 2'h0 & tempFraction[2] & (tempFraction[1] | tempFraction[0]) | _addOne_T_17; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 234:102]
  wire  _addOne_T_24 = tempFraction[2] | tempFraction[1] | tempFraction[0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 236:70]
  wire  _addOne_T_27 = roundingMode == 2'h1 & (tempFraction[2] | tempFraction[1] | tempFraction[0]) & resultSign; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 236:90]
  wire  _addOne_T_28 = _addOne_T_18 | _addOne_T_27; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 235:110]
  wire  _addOne_T_38 = roundingMode == 2'h2 & _addOne_T_24 & ~resultSign; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 237:90]
  wire  addOne = _addOne_T_28 | _addOne_T_38; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 236:106]
  wire [3:0] _GEN_16 = {{3'd0}, addOne}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 239:66]
  wire [4:0] roundedFraction = tempFraction[6:3] + _GEN_16; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 239:66]
  wire [3:0] resultFraction = roundedFraction[4] ? roundedFraction[4:1] : roundedFraction[3:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 241:28]
  wire [3:0] _finalExponent_T_7 = tempExponent + 4'h1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 245:20]
  wire [3:0] resultExponent = roundedFraction[4] | roundedFraction[3] & tempExponent == 4'h0 ? _finalExponent_T_7 :
    tempExponent; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 244:28]
  wire  _overflow_T_9 = tempExponent >= 4'hf & tempFraction[6:3] == 4'hf; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 250:42]
  wire  resultOverflow = resultExponent == 4'hf & resultFraction == 4'hf | _overflow_T_9; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 249:134]
  wire [3:0] _GEN_8 = enable ? resultExponent : 4'h0; // @[\\src\\main\\scala\\fpu8\\Add.scala 26:24 28:14 37:14]
  assign sign = enable & resultSign; // @[\\src\\main\\scala\\fpu8\\Add.scala 26:24 27:10 36:10]
  assign exponent = {{1'd0}, _GEN_8};
  assign fraction = enable ? resultFraction : 4'h0; // @[\\src\\main\\scala\\fpu8\\Add.scala 26:24 29:14 38:14]
  assign overflow = enable & resultOverflow; // @[\\src\\main\\scala\\fpu8\\Add.scala 26:24 30:14 39:14]
  assign is0 = enable & isResult0; // @[\\src\\main\\scala\\fpu8\\Add.scala 26:24 32:9 41:9]
  assign isNaN = enable & isResultNaN; // @[\\src\\main\\scala\\fpu8\\Add.scala 26:24 33:11 42:11]
endmodule
module Multiply(
  input        enable, // @[\\src\\main\\scala\\fpu8\\Multiply.scala 9:18]
  input  [7:0] a_data, // @[\\src\\main\\scala\\fpu8\\Multiply.scala 10:13]
  input  [7:0] b_data, // @[\\src\\main\\scala\\fpu8\\Multiply.scala 11:13]
  input  [1:0] roundingMode, // @[\\src\\main\\scala\\fpu8\\Multiply.scala 12:24]
  output       sign, // @[\\src\\main\\scala\\fpu8\\Multiply.scala 13:16]
  output [4:0] exponent, // @[\\src\\main\\scala\\fpu8\\Multiply.scala 14:20]
  output [3:0] fraction, // @[\\src\\main\\scala\\fpu8\\Multiply.scala 15:20]
  output       overflow, // @[\\src\\main\\scala\\fpu8\\Multiply.scala 16:20]
  output       is0, // @[\\src\\main\\scala\\fpu8\\Multiply.scala 18:15]
  output       isNaN // @[\\src\\main\\scala\\fpu8\\Multiply.scala 19:17]
);
  wire  _isResultNaN_T_1 = a_data[6:3] == 4'hf; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 35:41]
  wire  _isResultNaN_T_3 = a_data[2:0] == 3'h7; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 39:46]
  wire  _isResultNaN_T_4 = _isResultNaN_T_1 & _isResultNaN_T_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 41:30]
  wire  _isResultNaN_T_6 = b_data[6:3] == 4'hf; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 35:41]
  wire  _isResultNaN_T_8 = b_data[2:0] == 3'h7; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 39:46]
  wire  _isResultNaN_T_9 = _isResultNaN_T_6 & _isResultNaN_T_8; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 41:30]
  wire  isResultNaN = _isResultNaN_T_4 | _isResultNaN_T_9; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 441:37]
  wire  _isResult0_T_1 = a_data[6:3] == 4'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 33:39]
  wire  _isResult0_T_3 = a_data[2:0] == 3'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 37:44]
  wire  _isResult0_T_4 = _isResult0_T_1 & _isResult0_T_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 51:26]
  wire  _isResult0_T_13 = b_data[6:3] == 4'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 33:39]
  wire  _isResult0_T_15 = b_data[2:0] == 3'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 37:44]
  wire  _isResult0_T_16 = _isResult0_T_13 & _isResult0_T_15; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 51:26]
  wire  isResult0 = _isResult0_T_4 & ~_isResultNaN_T_9 | _isResult0_T_16 & ~_isResultNaN_T_4; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 449:62]
  wire  resultSign = a_data[7] ^ b_data[7]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 156:26]
  wire [5:0] _exponent_T_11 = {2'h0,a_data[6:3]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 162:16]
  wire [5:0] _exponent_T_13 = {2'h0,b_data[6:3]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 162:47]
  wire [5:0] _exponent_T_15 = _exponent_T_11 + _exponent_T_13; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 162:42]
  wire [5:0] _exponent_T_17 = _exponent_T_15 - 6'h6; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 162:74]
  wire [5:0] _exponent_T_25 = _exponent_T_15 - 6'h7; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 163:74]
  wire [5:0] _exponent_T_26 = _isResult0_T_1 ^ _isResult0_T_13 ? _exponent_T_17 : _exponent_T_25; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 161:14]
  wire [5:0] exponent_1 = _isResult0_T_1 & _isResult0_T_13 ? 6'h34 : _exponent_T_26; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 159:12]
  wire  _firstOperandFraction_T_2 = ~_isResult0_T_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 171:36]
  wire [3:0] firstOperandFraction = {_firstOperandFraction_T_2,a_data[2:0]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 171:35]
  wire  _secondOperandFraction_T_2 = ~_isResult0_T_13; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 172:37]
  wire [3:0] secondOperandFraction = {_secondOperandFraction_T_2,b_data[2:0]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 172:36]
  wire [3:0] product_partialProducts_compare = secondOperandFraction[0] ? 4'hf : 4'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 101:24]
  wire [3:0] product_partialProducts_0 = firstOperandFraction & product_partialProducts_compare; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:11]
  wire [3:0] product_partialProducts_compare_1 = secondOperandFraction[1] ? 4'hf : 4'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 101:24]
  wire [3:0] _product_partialProducts_T_1 = firstOperandFraction & product_partialProducts_compare_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:11]
  wire [4:0] product_partialProducts_1 = {_product_partialProducts_T_1, 1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:22]
  wire [3:0] product_partialProducts_compare_2 = secondOperandFraction[2] ? 4'hf : 4'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 101:24]
  wire [3:0] _product_partialProducts_T_2 = firstOperandFraction & product_partialProducts_compare_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:11]
  wire [5:0] product_partialProducts_2 = {_product_partialProducts_T_2, 2'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:22]
  wire [3:0] product_partialProducts_compare_3 = secondOperandFraction[3] ? 4'hf : 4'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 101:24]
  wire [3:0] _product_partialProducts_T_3 = firstOperandFraction & product_partialProducts_compare_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:11]
  wire [6:0] product_partialProducts_3 = {_product_partialProducts_T_3, 3'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:22]
  wire [4:0] _GEN_14 = {{1'd0}, product_partialProducts_0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 112:34]
  wire [5:0] _product_partialSums_T = _GEN_14 + product_partialProducts_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 112:34]
  wire [6:0] product_partialSums_0 = _product_partialSums_T + product_partialProducts_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 112:39]
  wire [7:0] product = product_partialSums_0 + product_partialProducts_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 109:15]
  wire [6:0] _leadingZeros_T_17 = {product[0],product[1],product[2],product[3],product[4],product[5],product[6]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 58:44]
  wire [2:0] _leadingZeros_T_25 = _leadingZeros_T_17[5] ? 3'h5 : 3'h6; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] _leadingZeros_T_26 = _leadingZeros_T_17[4] ? 3'h4 : _leadingZeros_T_25; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] _leadingZeros_T_27 = _leadingZeros_T_17[3] ? 3'h3 : _leadingZeros_T_26; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] _leadingZeros_T_28 = _leadingZeros_T_17[2] ? 3'h2 : _leadingZeros_T_27; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] _leadingZeros_T_29 = _leadingZeros_T_17[1] ? 3'h1 : _leadingZeros_T_28; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] shift = _leadingZeros_T_17[0] ? 3'h0 : _leadingZeros_T_29; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [7:0] _shiftedValue_T_3 = {product[6:0], 1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 63:23]
  wire [8:0] _shiftedValue_T_5 = {product[6:0], 2'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 63:23]
  wire [9:0] _shiftedValue_T_7 = {product[6:0], 3'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 63:23]
  wire [10:0] _shiftedValue_T_9 = {product[6:0], 4'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 63:23]
  wire [11:0] _shiftedValue_T_11 = {product[6:0], 5'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 63:23]
  wire [12:0] _shiftedValue_T_13 = {product[6:0], 6'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 63:23]
  wire [6:0] _shiftedValue_T_18 = 3'h1 == shift ? _shiftedValue_T_3[6:0] : product[6:0]; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [6:0] _shiftedValue_T_20 = 3'h2 == shift ? _shiftedValue_T_5[6:0] : _shiftedValue_T_18; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [6:0] _shiftedValue_T_22 = 3'h3 == shift ? _shiftedValue_T_7[6:0] : _shiftedValue_T_20; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [6:0] _shiftedValue_T_24 = 3'h4 == shift ? _shiftedValue_T_9[6:0] : _shiftedValue_T_22; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [6:0] _shiftedValue_T_26 = 3'h5 == shift ? _shiftedValue_T_11[6:0] : _shiftedValue_T_24; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [6:0] shiftedCalcValue = 3'h6 == shift ? _shiftedValue_T_13[6:0] : _shiftedValue_T_26; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [5:0] exponentShiftRight = 6'h0 - exponent_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 305:55]
  wire [5:0] exponentShiftLeft = exponent_1 - 6'h1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 308:35]
  wire  _T_2 = ~exponent_1[5]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 314:10]
  wire  _T_5 = ~exponent_1[5] & exponent_1[4:0] >= 5'hf; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 314:40]
  wire  _T_12 = _T_2 & exponent_1[4:0] < 5'hf; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 318:46]
  wire [4:0] _tempExponent_T_2 = exponent_1[4:0] + 5'h1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 320:38]
  wire [6:0] _tempFraction_T_3 = {product[7:2],|product[1:0]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 321:26]
  wire [4:0] _GEN_15 = {{2'd0}, shift}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 322:78]
  wire  _T_19 = _T_2 & exponent_1[4:0] > _GEN_15; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 322:46]
  wire [4:0] _tempExponent_T_5 = exponent_1[4:0] - _GEN_15; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 324:51]
  wire [6:0] _tempFraction_T_27 = 6'h0 == exponentShiftLeft ? product[6:0] : product[6:0]; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [6:0] _tempFraction_T_29 = 6'h1 == exponentShiftLeft ? _shiftedValue_T_3[6:0] : _tempFraction_T_27; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [6:0] _tempFraction_T_31 = 6'h2 == exponentShiftLeft ? _shiftedValue_T_5[6:0] : _tempFraction_T_29; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [6:0] _tempFraction_T_33 = 6'h3 == exponentShiftLeft ? _shiftedValue_T_7[6:0] : _tempFraction_T_31; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [6:0] _tempFraction_T_35 = 6'h4 == exponentShiftLeft ? _shiftedValue_T_9[6:0] : _tempFraction_T_33; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [6:0] _tempFraction_T_37 = 6'h5 == exponentShiftLeft ? _shiftedValue_T_11[6:0] : _tempFraction_T_35; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [6:0] _tempFraction_T_39 = 6'h6 == exponentShiftLeft ? _shiftedValue_T_13[6:0] : _tempFraction_T_37; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [6:0] _tempFraction_T_44 = _tempFraction_T_3 >> exponentShiftRight; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 336:110]
  wire [6:0] _GEN_0 = _T_2 & exponent_1[4:0] > 5'h0 ? _tempFraction_T_39 : _tempFraction_T_44; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 328:82 330:22 336:22]
  wire [4:0] _GEN_1 = _T_19 & shiftedCalcValue[6] ? _tempExponent_T_5 : 5'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 323:55 324:20 327:20]
  wire [6:0] _GEN_2 = _T_19 & shiftedCalcValue[6] ? shiftedCalcValue : _GEN_0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 323:55 325:20]
  wire [4:0] _GEN_3 = _T_12 & product[7] ? _tempExponent_T_2 : _GEN_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 319:54 320:20]
  wire [6:0] _GEN_4 = _T_12 & product[7] ? _tempFraction_T_3 : _GEN_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 319:54 321:20]
  wire [4:0] tempExponent = _T_5 & product[7] ? 5'hf : _GEN_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 315:54 316:20]
  wire [6:0] tempFraction = _T_5 & product[7] ? 7'h7f : _GEN_4; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 315:54 317:20]
  wire  _addOne_T_2 = roundingMode == 2'h0 & tempFraction[2]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 234:42]
  wire  _addOne_T_17 = _addOne_T_2 & ~tempFraction[1] & ~tempFraction[0] & tempFraction[3]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 235:90]
  wire  _addOne_T_18 = roundingMode == 2'h0 & tempFraction[2] & (tempFraction[1] | tempFraction[0]) | _addOne_T_17; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 234:102]
  wire  _addOne_T_24 = tempFraction[2] | tempFraction[1] | tempFraction[0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 236:70]
  wire  _addOne_T_27 = roundingMode == 2'h1 & (tempFraction[2] | tempFraction[1] | tempFraction[0]) & resultSign; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 236:90]
  wire  _addOne_T_28 = _addOne_T_18 | _addOne_T_27; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 235:110]
  wire  _addOne_T_38 = roundingMode == 2'h2 & _addOne_T_24 & ~resultSign; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 237:90]
  wire  addOne = _addOne_T_28 | _addOne_T_38; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 236:106]
  wire [3:0] _GEN_17 = {{3'd0}, addOne}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 239:66]
  wire [4:0] roundedFraction = tempFraction[6:3] + _GEN_17; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 239:66]
  wire [3:0] resultFraction = roundedFraction[4] ? roundedFraction[4:1] : roundedFraction[3:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 241:28]
  wire [4:0] _finalExponent_T_7 = tempExponent + 5'h1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 245:20]
  wire [4:0] resultExponent = roundedFraction[4] | roundedFraction[3] & tempExponent == 5'h0 ? _finalExponent_T_7 :
    tempExponent; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 244:28]
  wire  _overflow_T_9 = tempExponent >= 5'hf & tempFraction[6:3] == 4'hf; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 250:42]
  wire  resultOverflow = resultExponent > 5'hf | resultExponent[3:0] == 4'hf & resultFraction == 4'hf | _overflow_T_9; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 249:134]
  assign sign = enable & resultSign; // @[\\src\\main\\scala\\fpu8\\Multiply.scala 25:24 26:10 35:10]
  assign exponent = enable ? resultExponent : 5'h0; // @[\\src\\main\\scala\\fpu8\\Multiply.scala 25:24 27:14 36:14]
  assign fraction = enable ? resultFraction : 4'h0; // @[\\src\\main\\scala\\fpu8\\Multiply.scala 25:24 28:14 37:14]
  assign overflow = enable & resultOverflow; // @[\\src\\main\\scala\\fpu8\\Multiply.scala 25:24 29:14 38:14]
  assign is0 = enable & isResult0; // @[\\src\\main\\scala\\fpu8\\Multiply.scala 25:24 31:9 40:9]
  assign isNaN = enable & isResultNaN; // @[\\src\\main\\scala\\fpu8\\Multiply.scala 25:24 32:11 41:11]
endmodule
module Divide(
  input        enable, // @[\\src\\main\\scala\\fpu8\\Divide.scala 9:18]
  input  [7:0] a_data, // @[\\src\\main\\scala\\fpu8\\Divide.scala 10:13]
  input  [7:0] b_data, // @[\\src\\main\\scala\\fpu8\\Divide.scala 11:13]
  input  [1:0] roundingMode, // @[\\src\\main\\scala\\fpu8\\Divide.scala 12:24]
  output       sign, // @[\\src\\main\\scala\\fpu8\\Divide.scala 13:16]
  output [4:0] exponent, // @[\\src\\main\\scala\\fpu8\\Divide.scala 14:20]
  output [3:0] fraction, // @[\\src\\main\\scala\\fpu8\\Divide.scala 15:20]
  output       overflow, // @[\\src\\main\\scala\\fpu8\\Divide.scala 16:20]
  output       is0, // @[\\src\\main\\scala\\fpu8\\Divide.scala 18:15]
  output       isNaN // @[\\src\\main\\scala\\fpu8\\Divide.scala 19:17]
);
  wire  _isResultNaN_T_1 = a_data[6:3] == 4'hf; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 35:41]
  wire  _isResultNaN_T_3 = a_data[2:0] == 3'h7; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 39:46]
  wire  _isResultNaN_T_4 = _isResultNaN_T_1 & _isResultNaN_T_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 41:30]
  wire  _isResultNaN_T_6 = b_data[6:3] == 4'hf; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 35:41]
  wire  _isResultNaN_T_8 = b_data[2:0] == 3'h7; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 39:46]
  wire  _isResultNaN_T_9 = _isResultNaN_T_6 & _isResultNaN_T_8; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 41:30]
  wire  _isResultNaN_T_12 = b_data[6:3] == 4'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 33:39]
  wire  _isResultNaN_T_14 = b_data[2:0] == 3'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 37:44]
  wire  _isResultNaN_T_15 = _isResultNaN_T_12 & _isResultNaN_T_14; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 51:26]
  wire  isResultNaN = _isResultNaN_T_4 | _isResultNaN_T_9 | _isResultNaN_T_15; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 469:40]
  wire  _isResult0_T_1 = a_data[6:3] == 4'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 33:39]
  wire  _isResult0_T_3 = a_data[2:0] == 3'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 37:44]
  wire  _isResult0_T_4 = _isResult0_T_1 & _isResult0_T_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 51:26]
  wire  isResult0 = _isResult0_T_4 & ~_isResultNaN_T_15 & ~_isResultNaN_T_9; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 479:32]
  wire  resultSign = a_data[7] ^ b_data[7]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 178:26]
  wire [3:0] _tempDividendFraction_T_3 = {a_data[2:0],1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 180:10]
  wire [3:0] _tempDividendFraction_T_5 = {1'h1,a_data[2:0]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 181:10]
  wire [3:0] tempDividendFraction = _isResult0_T_1 ? _tempDividendFraction_T_3 : _tempDividendFraction_T_5; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 179:35]
  wire [3:0] _tempDivisorFraction_T_3 = {b_data[2:0],1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 184:10]
  wire [3:0] _tempDivisorFraction_T_5 = {1'h1,b_data[2:0]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 185:10]
  wire [3:0] tempDivisorFraction = _isResultNaN_T_12 ? _tempDivisorFraction_T_3 : _tempDivisorFraction_T_5; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 183:34]
  wire [5:0] _tempExponent_T_1 = {2'h0,a_data[6:3]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 187:27]
  wire [5:0] _tempExponent_T_3 = {2'h0,b_data[6:3]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 188:10]
  wire [5:0] _tempExponent_T_5 = _tempExponent_T_1 - _tempExponent_T_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 187:53]
  wire [5:0] tempExponent = _tempExponent_T_5 + 6'h7; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 188:37]
  wire [3:0] _leadingZeros_T_8 = {tempDividendFraction[0],tempDividendFraction[1],tempDividendFraction[2],
    tempDividendFraction[3]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 58:44]
  wire [1:0] _leadingZeros_T_13 = _leadingZeros_T_8[2] ? 2'h2 : 2'h3; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [1:0] _leadingZeros_T_14 = _leadingZeros_T_8[1] ? 2'h1 : _leadingZeros_T_13; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [1:0] dividendShift = _leadingZeros_T_8[0] ? 2'h0 : _leadingZeros_T_14; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _shiftedValue_T_3 = {tempDividendFraction, 1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 63:23]
  wire [5:0] _shiftedValue_T_5 = {tempDividendFraction, 2'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 63:23]
  wire [6:0] _shiftedValue_T_7 = {tempDividendFraction, 3'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 63:23]
  wire [3:0] _shiftedValue_T_10 = 2'h1 == dividendShift ? _shiftedValue_T_3[3:0] : tempDividendFraction; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [3:0] _shiftedValue_T_12 = 2'h2 == dividendShift ? _shiftedValue_T_5[3:0] : _shiftedValue_T_10; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [3:0] dividendFraction = 2'h3 == dividendShift ? _shiftedValue_T_7[3:0] : _shiftedValue_T_12; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [3:0] _leadingZeros_T_24 = {tempDivisorFraction[0],tempDivisorFraction[1],tempDivisorFraction[2],
    tempDivisorFraction[3]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 58:44]
  wire [1:0] _leadingZeros_T_29 = _leadingZeros_T_24[2] ? 2'h2 : 2'h3; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [1:0] _leadingZeros_T_30 = _leadingZeros_T_24[1] ? 2'h1 : _leadingZeros_T_29; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [1:0] divisorShift = _leadingZeros_T_24[0] ? 2'h0 : _leadingZeros_T_30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _shiftedValue_T_18 = {tempDivisorFraction, 1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 63:23]
  wire [5:0] _shiftedValue_T_20 = {tempDivisorFraction, 2'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 63:23]
  wire [6:0] _shiftedValue_T_22 = {tempDivisorFraction, 3'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 63:23]
  wire [3:0] _shiftedValue_T_25 = 2'h1 == divisorShift ? _shiftedValue_T_18[3:0] : tempDivisorFraction; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [3:0] _shiftedValue_T_27 = 2'h2 == divisorShift ? _shiftedValue_T_20[3:0] : _shiftedValue_T_25; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [3:0] divisorFraction = 2'h3 == divisorShift ? _shiftedValue_T_22[3:0] : _shiftedValue_T_27; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [5:0] _GEN_22 = {{4'd0}, dividendShift}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 195:33]
  wire [5:0] _exponent_T_1 = tempExponent - _GEN_22; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 195:33]
  wire [5:0] _GEN_23 = {{4'd0}, divisorShift}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 195:49]
  wire [5:0] exponent_1 = _exponent_T_1 + _GEN_23; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 195:49]
  wire [3:0] _GEN_1 = 3'h1 == divisorFraction[2:0] ? 4'hc : 4'he; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 203:{24,24}]
  wire [3:0] _GEN_2 = 3'h2 == divisorFraction[2:0] ? 4'ha : _GEN_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 203:{24,24}]
  wire [3:0] _GEN_3 = 3'h3 == divisorFraction[2:0] ? 4'h8 : _GEN_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 203:{24,24}]
  wire [3:0] _GEN_4 = 3'h4 == divisorFraction[2:0] ? 4'h6 : _GEN_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 203:{24,24}]
  wire [3:0] _GEN_5 = 3'h5 == divisorFraction[2:0] ? 4'h4 : _GEN_4; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 203:{24,24}]
  wire [3:0] _GEN_6 = 3'h6 == divisorFraction[2:0] ? 4'h2 : _GEN_5; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 203:{24,24}]
  wire [3:0] _GEN_7 = 3'h7 == divisorFraction[2:0] ? 4'h0 : _GEN_6; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 203:{24,24}]
  wire [5:0] quotient_initGuess = {2'h1,_GEN_7}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 203:24]
  wire [5:0] quotient_secondGuess_firstStep_partialProducts_compare = divisorFraction[0] ? 6'h3f : 6'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 101:24]
  wire [5:0] quotient_secondGuess_firstStep_partialProducts_0 = quotient_initGuess &
    quotient_secondGuess_firstStep_partialProducts_compare; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:11]
  wire [5:0] quotient_secondGuess_firstStep_partialProducts_compare_1 = divisorFraction[1] ? 6'h3f : 6'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 101:24]
  wire [5:0] _quotient_secondGuess_firstStep_partialProducts_T_1 = quotient_initGuess &
    quotient_secondGuess_firstStep_partialProducts_compare_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:11]
  wire [6:0] quotient_secondGuess_firstStep_partialProducts_1 = {_quotient_secondGuess_firstStep_partialProducts_T_1
    , 1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:22]
  wire [5:0] quotient_secondGuess_firstStep_partialProducts_compare_2 = divisorFraction[2] ? 6'h3f : 6'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 101:24]
  wire [5:0] _quotient_secondGuess_firstStep_partialProducts_T_2 = quotient_initGuess &
    quotient_secondGuess_firstStep_partialProducts_compare_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:11]
  wire [7:0] quotient_secondGuess_firstStep_partialProducts_2 = {_quotient_secondGuess_firstStep_partialProducts_T_2
    , 2'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:22]
  wire [5:0] quotient_secondGuess_firstStep_partialProducts_compare_3 = divisorFraction[3] ? 6'h3f : 6'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 101:24]
  wire [5:0] _quotient_secondGuess_firstStep_partialProducts_T_3 = quotient_initGuess &
    quotient_secondGuess_firstStep_partialProducts_compare_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:11]
  wire [8:0] quotient_secondGuess_firstStep_partialProducts_3 = {_quotient_secondGuess_firstStep_partialProducts_T_3
    , 3'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:22]
  wire [6:0] _GEN_24 = {{1'd0}, quotient_secondGuess_firstStep_partialProducts_0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 112:34]
  wire [7:0] _quotient_secondGuess_firstStep_partialSums_T = _GEN_24 + quotient_secondGuess_firstStep_partialProducts_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 112:34]
  wire [8:0] quotient_secondGuess_firstStep_partialSums_0 = _quotient_secondGuess_firstStep_partialSums_T +
    quotient_secondGuess_firstStep_partialProducts_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 112:39]
  wire [9:0] quotient_secondGuess_firstStep = quotient_secondGuess_firstStep_partialSums_0 +
    quotient_secondGuess_firstStep_partialProducts_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 109:15]
  wire  _quotient_secondGuess_firstStepRnd_roundedValue_T_4 = quotient_secondGuess_firstStep[2] & |
    quotient_secondGuess_firstStep[1:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 77:59]
  wire [5:0] _GEN_25 = {{5'd0}, _quotient_secondGuess_firstStepRnd_roundedValue_T_4}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 77:35]
  wire [6:0] quotient_secondGuess_firstStepRnd = quotient_secondGuess_firstStep[8:3] + _GEN_25; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 77:35]
  wire [5:0] _quotient_secondGuess_secondStep_T_1 = ~quotient_secondGuess_firstStepRnd[5:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 214:25]
  wire [5:0] quotient_secondGuess_secondStep = _quotient_secondGuess_secondStep_T_1 + 6'h1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 214:70]
  wire [5:0] quotient_secondGuess_finalStep_partialProducts_compare = quotient_secondGuess_secondStep[0] ? 6'h3f : 6'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 101:24]
  wire [5:0] quotient_secondGuess_finalStep_partialProducts_0 = quotient_initGuess &
    quotient_secondGuess_finalStep_partialProducts_compare; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:11]
  wire [5:0] quotient_secondGuess_finalStep_partialProducts_compare_1 = quotient_secondGuess_secondStep[1] ? 6'h3f : 6'h0
    ; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 101:24]
  wire [5:0] _quotient_secondGuess_finalStep_partialProducts_T_1 = quotient_initGuess &
    quotient_secondGuess_finalStep_partialProducts_compare_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:11]
  wire [6:0] quotient_secondGuess_finalStep_partialProducts_1 = {_quotient_secondGuess_finalStep_partialProducts_T_1
    , 1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:22]
  wire [5:0] quotient_secondGuess_finalStep_partialProducts_compare_2 = quotient_secondGuess_secondStep[2] ? 6'h3f : 6'h0
    ; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 101:24]
  wire [5:0] _quotient_secondGuess_finalStep_partialProducts_T_2 = quotient_initGuess &
    quotient_secondGuess_finalStep_partialProducts_compare_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:11]
  wire [7:0] quotient_secondGuess_finalStep_partialProducts_2 = {_quotient_secondGuess_finalStep_partialProducts_T_2
    , 2'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:22]
  wire [5:0] quotient_secondGuess_finalStep_partialProducts_compare_3 = quotient_secondGuess_secondStep[3] ? 6'h3f : 6'h0
    ; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 101:24]
  wire [5:0] _quotient_secondGuess_finalStep_partialProducts_T_3 = quotient_initGuess &
    quotient_secondGuess_finalStep_partialProducts_compare_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:11]
  wire [8:0] quotient_secondGuess_finalStep_partialProducts_3 = {_quotient_secondGuess_finalStep_partialProducts_T_3
    , 3'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:22]
  wire [5:0] quotient_secondGuess_finalStep_partialProducts_compare_4 = quotient_secondGuess_secondStep[4] ? 6'h3f : 6'h0
    ; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 101:24]
  wire [5:0] _quotient_secondGuess_finalStep_partialProducts_T_4 = quotient_initGuess &
    quotient_secondGuess_finalStep_partialProducts_compare_4; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:11]
  wire [9:0] quotient_secondGuess_finalStep_partialProducts_4 = {_quotient_secondGuess_finalStep_partialProducts_T_4
    , 4'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:22]
  wire [5:0] quotient_secondGuess_finalStep_partialProducts_compare_5 = quotient_secondGuess_secondStep[5] ? 6'h3f : 6'h0
    ; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 101:24]
  wire [5:0] _quotient_secondGuess_finalStep_partialProducts_T_5 = quotient_initGuess &
    quotient_secondGuess_finalStep_partialProducts_compare_5; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:11]
  wire [10:0] quotient_secondGuess_finalStep_partialProducts_5 = {_quotient_secondGuess_finalStep_partialProducts_T_5
    , 5'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:22]
  wire [6:0] _GEN_26 = {{1'd0}, quotient_secondGuess_finalStep_partialProducts_0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 112:34]
  wire [7:0] _quotient_secondGuess_finalStep_partialSums_T = _GEN_26 + quotient_secondGuess_finalStep_partialProducts_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 112:34]
  wire [8:0] quotient_secondGuess_finalStep_partialSums_0 = _quotient_secondGuess_finalStep_partialSums_T +
    quotient_secondGuess_finalStep_partialProducts_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 112:39]
  wire [9:0] _GEN_27 = {{1'd0}, quotient_secondGuess_finalStep_partialProducts_3}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 112:34]
  wire [10:0] _quotient_secondGuess_finalStep_partialSums_T_1 = _GEN_27 +
    quotient_secondGuess_finalStep_partialProducts_4; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 112:34]
  wire [11:0] quotient_secondGuess_finalStep_partialSums_1 = _quotient_secondGuess_finalStep_partialSums_T_1 +
    quotient_secondGuess_finalStep_partialProducts_5; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 112:39]
  wire [11:0] _GEN_28 = {{3'd0}, quotient_secondGuess_finalStep_partialSums_0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 109:15]
  wire [12:0] _quotient_secondGuess_finalStep_T = _GEN_28 + quotient_secondGuess_finalStep_partialSums_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 109:15]
  wire [11:0] quotient_secondGuess_finalStep = _quotient_secondGuess_finalStep_T[11:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 218:27 219:17]
  wire  _quotient_secondGuess_res_roundedValue_T_4 = quotient_secondGuess_finalStep[4] & |quotient_secondGuess_finalStep
    [3:2]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 77:59]
  wire [5:0] _GEN_29 = {{5'd0}, _quotient_secondGuess_res_roundedValue_T_4}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 77:35]
  wire [6:0] quotient_secondGuess = quotient_secondGuess_finalStep[10:5] + _GEN_29; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 77:35]
  wire [5:0] quotient_finalGuess_firstStep_partialProducts_0 = quotient_secondGuess[5:0] &
    quotient_secondGuess_firstStep_partialProducts_compare; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:11]
  wire [5:0] _quotient_finalGuess_firstStep_partialProducts_T_1 = quotient_secondGuess[5:0] &
    quotient_secondGuess_firstStep_partialProducts_compare_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:11]
  wire [6:0] quotient_finalGuess_firstStep_partialProducts_1 = {_quotient_finalGuess_firstStep_partialProducts_T_1
    , 1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:22]
  wire [5:0] _quotient_finalGuess_firstStep_partialProducts_T_2 = quotient_secondGuess[5:0] &
    quotient_secondGuess_firstStep_partialProducts_compare_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:11]
  wire [7:0] quotient_finalGuess_firstStep_partialProducts_2 = {_quotient_finalGuess_firstStep_partialProducts_T_2
    , 2'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:22]
  wire [5:0] _quotient_finalGuess_firstStep_partialProducts_T_3 = quotient_secondGuess[5:0] &
    quotient_secondGuess_firstStep_partialProducts_compare_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:11]
  wire [8:0] quotient_finalGuess_firstStep_partialProducts_3 = {_quotient_finalGuess_firstStep_partialProducts_T_3
    , 3'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:22]
  wire [6:0] _GEN_30 = {{1'd0}, quotient_finalGuess_firstStep_partialProducts_0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 112:34]
  wire [7:0] _quotient_finalGuess_firstStep_partialSums_T = _GEN_30 + quotient_finalGuess_firstStep_partialProducts_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 112:34]
  wire [8:0] quotient_finalGuess_firstStep_partialSums_0 = _quotient_finalGuess_firstStep_partialSums_T +
    quotient_finalGuess_firstStep_partialProducts_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 112:39]
  wire [9:0] quotient_finalGuess_firstStep = quotient_finalGuess_firstStep_partialSums_0 +
    quotient_finalGuess_firstStep_partialProducts_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 109:15]
  wire  _quotient_finalGuess_firstStepRnd_roundedValue_T_4 = quotient_finalGuess_firstStep[2] & |
    quotient_finalGuess_firstStep[1:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 77:59]
  wire [5:0] _GEN_31 = {{5'd0}, _quotient_finalGuess_firstStepRnd_roundedValue_T_4}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 77:35]
  wire [6:0] quotient_finalGuess_firstStepRnd = quotient_finalGuess_firstStep[8:3] + _GEN_31; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 77:35]
  wire [5:0] _quotient_finalGuess_secondStep_T_1 = ~quotient_finalGuess_firstStepRnd[5:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 214:25]
  wire [5:0] quotient_finalGuess_secondStep = _quotient_finalGuess_secondStep_T_1 + 6'h1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 214:70]
  wire [5:0] quotient_finalGuess_finalStep_partialProducts_compare = quotient_finalGuess_secondStep[0] ? 6'h3f : 6'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 101:24]
  wire [5:0] quotient_finalGuess_finalStep_partialProducts_0 = quotient_secondGuess[5:0] &
    quotient_finalGuess_finalStep_partialProducts_compare; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:11]
  wire [5:0] quotient_finalGuess_finalStep_partialProducts_compare_1 = quotient_finalGuess_secondStep[1] ? 6'h3f : 6'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 101:24]
  wire [5:0] _quotient_finalGuess_finalStep_partialProducts_T_1 = quotient_secondGuess[5:0] &
    quotient_finalGuess_finalStep_partialProducts_compare_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:11]
  wire [6:0] quotient_finalGuess_finalStep_partialProducts_1 = {_quotient_finalGuess_finalStep_partialProducts_T_1
    , 1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:22]
  wire [5:0] quotient_finalGuess_finalStep_partialProducts_compare_2 = quotient_finalGuess_secondStep[2] ? 6'h3f : 6'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 101:24]
  wire [5:0] _quotient_finalGuess_finalStep_partialProducts_T_2 = quotient_secondGuess[5:0] &
    quotient_finalGuess_finalStep_partialProducts_compare_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:11]
  wire [7:0] quotient_finalGuess_finalStep_partialProducts_2 = {_quotient_finalGuess_finalStep_partialProducts_T_2
    , 2'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:22]
  wire [5:0] quotient_finalGuess_finalStep_partialProducts_compare_3 = quotient_finalGuess_secondStep[3] ? 6'h3f : 6'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 101:24]
  wire [5:0] _quotient_finalGuess_finalStep_partialProducts_T_3 = quotient_secondGuess[5:0] &
    quotient_finalGuess_finalStep_partialProducts_compare_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:11]
  wire [8:0] quotient_finalGuess_finalStep_partialProducts_3 = {_quotient_finalGuess_finalStep_partialProducts_T_3
    , 3'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:22]
  wire [5:0] quotient_finalGuess_finalStep_partialProducts_compare_4 = quotient_finalGuess_secondStep[4] ? 6'h3f : 6'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 101:24]
  wire [5:0] _quotient_finalGuess_finalStep_partialProducts_T_4 = quotient_secondGuess[5:0] &
    quotient_finalGuess_finalStep_partialProducts_compare_4; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:11]
  wire [9:0] quotient_finalGuess_finalStep_partialProducts_4 = {_quotient_finalGuess_finalStep_partialProducts_T_4
    , 4'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:22]
  wire [5:0] quotient_finalGuess_finalStep_partialProducts_compare_5 = quotient_finalGuess_secondStep[5] ? 6'h3f : 6'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 101:24]
  wire [5:0] _quotient_finalGuess_finalStep_partialProducts_T_5 = quotient_secondGuess[5:0] &
    quotient_finalGuess_finalStep_partialProducts_compare_5; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:11]
  wire [10:0] quotient_finalGuess_finalStep_partialProducts_5 = {_quotient_finalGuess_finalStep_partialProducts_T_5
    , 5'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:22]
  wire [6:0] _GEN_32 = {{1'd0}, quotient_finalGuess_finalStep_partialProducts_0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 112:34]
  wire [7:0] _quotient_finalGuess_finalStep_partialSums_T = _GEN_32 + quotient_finalGuess_finalStep_partialProducts_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 112:34]
  wire [8:0] quotient_finalGuess_finalStep_partialSums_0 = _quotient_finalGuess_finalStep_partialSums_T +
    quotient_finalGuess_finalStep_partialProducts_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 112:39]
  wire [9:0] _GEN_33 = {{1'd0}, quotient_finalGuess_finalStep_partialProducts_3}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 112:34]
  wire [10:0] _quotient_finalGuess_finalStep_partialSums_T_1 = _GEN_33 + quotient_finalGuess_finalStep_partialProducts_4
    ; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 112:34]
  wire [11:0] quotient_finalGuess_finalStep_partialSums_1 = _quotient_finalGuess_finalStep_partialSums_T_1 +
    quotient_finalGuess_finalStep_partialProducts_5; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 112:39]
  wire [11:0] _GEN_34 = {{3'd0}, quotient_finalGuess_finalStep_partialSums_0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 109:15]
  wire [12:0] _quotient_finalGuess_finalStep_T = _GEN_34 + quotient_finalGuess_finalStep_partialSums_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 109:15]
  wire [11:0] quotient_finalGuess_finalStep = _quotient_finalGuess_finalStep_T[11:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 218:27 219:17]
  wire  _quotient_finalGuess_res_roundedValue_T_4 = quotient_finalGuess_finalStep[4] & |quotient_finalGuess_finalStep[3:
    2]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 77:59]
  wire [5:0] _GEN_35 = {{5'd0}, _quotient_finalGuess_res_roundedValue_T_4}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 77:35]
  wire [6:0] quotient_finalGuess = quotient_finalGuess_finalStep[10:5] + _GEN_35; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 77:35]
  wire [5:0] quotient_partialProducts_compare = dividendFraction[0] ? 6'h3f : 6'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 101:24]
  wire [5:0] quotient_partialProducts_0 = quotient_finalGuess[5:0] & quotient_partialProducts_compare; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:11]
  wire [5:0] quotient_partialProducts_compare_1 = dividendFraction[1] ? 6'h3f : 6'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 101:24]
  wire [5:0] _quotient_partialProducts_T_1 = quotient_finalGuess[5:0] & quotient_partialProducts_compare_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:11]
  wire [6:0] quotient_partialProducts_1 = {_quotient_partialProducts_T_1, 1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:22]
  wire [5:0] quotient_partialProducts_compare_2 = dividendFraction[2] ? 6'h3f : 6'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 101:24]
  wire [5:0] _quotient_partialProducts_T_2 = quotient_finalGuess[5:0] & quotient_partialProducts_compare_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:11]
  wire [7:0] quotient_partialProducts_2 = {_quotient_partialProducts_T_2, 2'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:22]
  wire [5:0] quotient_partialProducts_compare_3 = dividendFraction[3] ? 6'h3f : 6'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 101:24]
  wire [5:0] _quotient_partialProducts_T_3 = quotient_finalGuess[5:0] & quotient_partialProducts_compare_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:11]
  wire [8:0] quotient_partialProducts_3 = {_quotient_partialProducts_T_3, 3'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:22]
  wire [6:0] _GEN_36 = {{1'd0}, quotient_partialProducts_0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 112:34]
  wire [7:0] _quotient_partialSums_T = _GEN_36 + quotient_partialProducts_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 112:34]
  wire [8:0] quotient_partialSums_0 = _quotient_partialSums_T + quotient_partialProducts_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 112:39]
  wire [9:0] quotient = quotient_partialSums_0 + quotient_partialProducts_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 109:15]
  wire [7:0] _GEN_37 = {{4'd0}, quotient[7:4]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 58:44]
  wire [7:0] _leadingZeros_T_36 = _GEN_37 & 8'hf; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 58:44]
  wire [7:0] _leadingZeros_T_38 = {quotient[3:0], 4'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 58:44]
  wire [7:0] _leadingZeros_T_40 = _leadingZeros_T_38 & 8'hf0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 58:44]
  wire [7:0] _leadingZeros_T_41 = _leadingZeros_T_36 | _leadingZeros_T_40; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 58:44]
  wire [7:0] _GEN_38 = {{2'd0}, _leadingZeros_T_41[7:2]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 58:44]
  wire [7:0] _leadingZeros_T_46 = _GEN_38 & 8'h33; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 58:44]
  wire [7:0] _leadingZeros_T_48 = {_leadingZeros_T_41[5:0], 2'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 58:44]
  wire [7:0] _leadingZeros_T_50 = _leadingZeros_T_48 & 8'hcc; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 58:44]
  wire [7:0] _leadingZeros_T_51 = _leadingZeros_T_46 | _leadingZeros_T_50; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 58:44]
  wire [7:0] _GEN_39 = {{1'd0}, _leadingZeros_T_51[7:1]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 58:44]
  wire [7:0] _leadingZeros_T_56 = _GEN_39 & 8'h55; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 58:44]
  wire [7:0] _leadingZeros_T_58 = {_leadingZeros_T_51[6:0], 1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 58:44]
  wire [7:0] _leadingZeros_T_60 = _leadingZeros_T_58 & 8'haa; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 58:44]
  wire [7:0] _leadingZeros_T_61 = _leadingZeros_T_56 | _leadingZeros_T_60; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 58:44]
  wire [8:0] _leadingZeros_T_63 = {_leadingZeros_T_61,quotient[8]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 58:44]
  wire [3:0] _leadingZeros_T_73 = _leadingZeros_T_63[7] ? 4'h7 : 4'h8; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _leadingZeros_T_74 = _leadingZeros_T_63[6] ? 4'h6 : _leadingZeros_T_73; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _leadingZeros_T_75 = _leadingZeros_T_63[5] ? 4'h5 : _leadingZeros_T_74; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _leadingZeros_T_76 = _leadingZeros_T_63[4] ? 4'h4 : _leadingZeros_T_75; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _leadingZeros_T_77 = _leadingZeros_T_63[3] ? 4'h3 : _leadingZeros_T_76; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _leadingZeros_T_78 = _leadingZeros_T_63[2] ? 4'h2 : _leadingZeros_T_77; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _leadingZeros_T_79 = _leadingZeros_T_63[1] ? 4'h1 : _leadingZeros_T_78; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] shift = _leadingZeros_T_63[0] ? 4'h0 : _leadingZeros_T_79; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [9:0] _shiftedValue_T_33 = {quotient[8:0], 1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 63:23]
  wire [10:0] _shiftedValue_T_35 = {quotient[8:0], 2'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 63:23]
  wire [11:0] _shiftedValue_T_37 = {quotient[8:0], 3'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 63:23]
  wire [12:0] _shiftedValue_T_39 = {quotient[8:0], 4'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 63:23]
  wire [13:0] _shiftedValue_T_41 = {quotient[8:0], 5'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 63:23]
  wire [14:0] _shiftedValue_T_43 = {quotient[8:0], 6'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 63:23]
  wire [15:0] _shiftedValue_T_45 = {quotient[8:0], 7'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 63:23]
  wire [16:0] _shiftedValue_T_47 = {quotient[8:0], 8'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 63:23]
  wire [8:0] _shiftedValue_T_52 = 4'h1 == shift ? _shiftedValue_T_33[8:0] : quotient[8:0]; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [8:0] _shiftedValue_T_54 = 4'h2 == shift ? _shiftedValue_T_35[8:0] : _shiftedValue_T_52; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [8:0] _shiftedValue_T_56 = 4'h3 == shift ? _shiftedValue_T_37[8:0] : _shiftedValue_T_54; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [8:0] _shiftedValue_T_58 = 4'h4 == shift ? _shiftedValue_T_39[8:0] : _shiftedValue_T_56; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [8:0] _shiftedValue_T_60 = 4'h5 == shift ? _shiftedValue_T_41[8:0] : _shiftedValue_T_58; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [8:0] _shiftedValue_T_62 = 4'h6 == shift ? _shiftedValue_T_43[8:0] : _shiftedValue_T_60; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [8:0] _shiftedValue_T_64 = 4'h7 == shift ? _shiftedValue_T_45[8:0] : _shiftedValue_T_62; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [8:0] shiftedCalcValue = 4'h8 == shift ? _shiftedValue_T_47[8:0] : _shiftedValue_T_64; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [5:0] exponentShiftRight = 6'h0 - exponent_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 352:55]
  wire [5:0] exponentShiftLeft = exponent_1 - 6'h1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 355:35]
  wire  _T_2 = ~exponent_1[5]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 363:10]
  wire  _T_5 = ~exponent_1[5] & exponent_1[4:0] >= 5'hf; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 363:40]
  wire  _T_12 = _T_2 & exponent_1[4:0] < 5'hf; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 367:46]
  wire [4:0] _tempExponent_T_9 = exponent_1[4:0] + 5'h1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 369:51]
  wire  _tempFraction_T_2 = &quotient[1:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 373:59]
  wire [6:0] _GEN_40 = {{6'd0}, _tempFraction_T_2}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 372:81]
  wire [6:0] _tempFraction_T_4 = quotient[8:2] + _GEN_40; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 372:81]
  wire [4:0] _GEN_41 = {{1'd0}, shift}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 377:78]
  wire  _T_19 = _T_2 & exponent_1[4:0] > _GEN_41; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 377:46]
  wire [4:0] _tempExponent_T_12 = exponent_1[4:0] - _GEN_41; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 379:51]
  wire  _tempFraction_T_7 = &shiftedCalcValue[1:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 383:60]
  wire [6:0] _GEN_43 = {{6'd0}, _tempFraction_T_7}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 382:82]
  wire [6:0] _tempFraction_T_9 = shiftedCalcValue[8:2] + _GEN_43; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 382:82]
  wire [69:0] _GEN_0 = {{63'd0}, _tempFraction_T_4}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 393:74]
  wire [69:0] _tempFraction_T_15 = _GEN_0 << exponentShiftLeft; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 393:74]
  wire  _tempFraction_T_18 = &quotient[2:1]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 399:125]
  wire [6:0] _GEN_45 = {{6'd0}, _tempFraction_T_18}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 398:118]
  wire [6:0] _tempFraction_T_20 = quotient[9:3] + _GEN_45; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 398:118]
  wire [6:0] _tempFraction_T_21 = _tempFraction_T_20 >> exponentShiftRight; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 399:138]
  wire [69:0] _GEN_8 = _T_2 & exponent_1[4:0] > 5'h0 ? _tempFraction_T_15 : {{63'd0}, _tempFraction_T_21}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 389:82 390:22 398:22]
  wire [4:0] _GEN_9 = _T_19 & shiftedCalcValue[8] ? _tempExponent_T_12 : 5'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 378:55 379:20 388:20]
  wire [69:0] _GEN_10 = _T_19 & shiftedCalcValue[8] ? {{63'd0}, _tempFraction_T_9} : _GEN_8; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 378:55 380:20]
  wire [4:0] _GEN_11 = _T_12 & quotient[9] ? _tempExponent_T_9 : _GEN_9; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 368:54 369:20]
  wire [69:0] _GEN_12 = _T_12 & quotient[9] ? {{63'd0}, _tempFraction_T_4} : _GEN_10; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 368:54 370:20]
  wire [4:0] tempExponent_1 = _T_5 & quotient[9] ? 5'hf : _GEN_11; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 364:54 365:20]
  wire [69:0] _GEN_14 = _T_5 & quotient[9] ? 70'hff : _GEN_12; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 364:54 366:20]
  wire [7:0] tempFraction = _GEN_14[7:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 359:28]
  wire  _addOne_T_2 = roundingMode == 2'h0 & tempFraction[2]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 234:42]
  wire  _addOne_T_17 = _addOne_T_2 & ~tempFraction[1] & ~tempFraction[0] & tempFraction[3]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 235:90]
  wire  _addOne_T_18 = roundingMode == 2'h0 & tempFraction[2] & (tempFraction[1] | tempFraction[0]) | _addOne_T_17; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 234:102]
  wire  _addOne_T_24 = tempFraction[2] | tempFraction[1] | tempFraction[0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 236:70]
  wire  _addOne_T_27 = roundingMode == 2'h1 & (tempFraction[2] | tempFraction[1] | tempFraction[0]) & resultSign; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 236:90]
  wire  _addOne_T_28 = _addOne_T_18 | _addOne_T_27; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 235:110]
  wire  _addOne_T_38 = roundingMode == 2'h2 & _addOne_T_24 & ~resultSign; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 237:90]
  wire  addOne = _addOne_T_28 | _addOne_T_38; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 236:106]
  wire [3:0] _GEN_46 = {{3'd0}, addOne}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 239:66]
  wire [4:0] roundedFraction = tempFraction[6:3] + _GEN_46; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 239:66]
  wire [3:0] resultFraction = roundedFraction[4] ? roundedFraction[4:1] : roundedFraction[3:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 241:28]
  wire [4:0] _finalExponent_T_7 = tempExponent_1 + 5'h1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 245:20]
  wire [4:0] resultExponent = roundedFraction[4] | roundedFraction[3] & tempExponent_1 == 5'h0 ? _finalExponent_T_7 :
    tempExponent_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 244:28]
  wire  _overflow_T_9 = tempExponent_1 >= 5'hf & tempFraction[6:3] == 4'hf; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 250:42]
  wire  resultOverflow = resultExponent > 5'hf | resultExponent[3:0] == 4'hf & resultFraction == 4'hf | _overflow_T_9; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 249:134]
  assign sign = enable & resultSign; // @[\\src\\main\\scala\\fpu8\\Divide.scala 25:24 26:10 35:10]
  assign exponent = enable ? resultExponent : 5'h0; // @[\\src\\main\\scala\\fpu8\\Divide.scala 25:24 27:14 36:14]
  assign fraction = enable ? resultFraction : 4'h0; // @[\\src\\main\\scala\\fpu8\\Divide.scala 25:24 28:14 37:14]
  assign overflow = enable & resultOverflow; // @[\\src\\main\\scala\\fpu8\\Divide.scala 25:24 29:14 38:14]
  assign is0 = enable & isResult0; // @[\\src\\main\\scala\\fpu8\\Divide.scala 25:24 31:9 40:9]
  assign isNaN = enable & isResultNaN; // @[\\src\\main\\scala\\fpu8\\Divide.scala 25:24 32:11 41:11]
endmodule
module Compare(
  input        enable, // @[\\src\\main\\scala\\fpu8\\Compare.scala 6:18]
  input  [2:0] compareMode, // @[\\src\\main\\scala\\fpu8\\Compare.scala 7:23]
  input  [7:0] a_data, // @[\\src\\main\\scala\\fpu8\\Compare.scala 8:13]
  input  [7:0] b_data, // @[\\src\\main\\scala\\fpu8\\Compare.scala 9:13]
  output [7:0] z // @[\\src\\main\\scala\\fpu8\\Compare.scala 10:13]
);
  wire  _z_isResultNaN_T_1 = a_data[6:3] == 4'hf; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 35:41]
  wire  _z_isResultNaN_T_3 = a_data[2:0] == 3'h7; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 39:46]
  wire  _z_isResultNaN_T_4 = _z_isResultNaN_T_1 & _z_isResultNaN_T_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 41:30]
  wire  _z_isResultNaN_T_6 = b_data[6:3] == 4'hf; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 35:41]
  wire  _z_isResultNaN_T_8 = b_data[2:0] == 3'h7; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 39:46]
  wire  _z_isResultNaN_T_9 = _z_isResultNaN_T_6 & _z_isResultNaN_T_8; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 41:30]
  wire  z_isResultNaN = _z_isResultNaN_T_4 | _z_isResultNaN_T_9; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 498:34]
  wire  _z_T_7 = a_data[6:0] > b_data[6:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 29:77]
  wire  _z_T_11 = ~a_data[7]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 506:102]
  wire  _z_T_15 = ~_z_T_7; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 506:113]
  wire [7:0] _GEN_0 = a_data[7] > b_data[7] | a_data[7] & _z_T_7 | ~a_data[7] & ~_z_T_7 ? 8'h38 : 8'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 506:138 508:14 510:14]
  wire [7:0] z_result = z_isResultNaN ? 8'h7f : _GEN_0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 501:22 502:14]
  wire [7:0] _GEN_2 = a_data[7] < b_data[7] | a_data[7] & _z_T_15 | _z_T_11 & _z_T_7 ? 8'h38 : 8'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 527:139 529:14 531:14]
  wire [7:0] z_result_1 = z_isResultNaN ? 8'h7f : _GEN_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 522:22 523:14]
  wire [7:0] _GEN_4 = a_data == b_data ? 8'h38 : 8'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 548:42 550:14 552:14]
  wire [7:0] z_result_2 = z_isResultNaN ? 8'h7f : _GEN_4; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 543:23 544:14]
  wire [7:0] _z_result_T_26 = z_result ^ z_result_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 570:32]
  wire [7:0] z_result_3 = z_isResultNaN ? 8'h7f : _z_result_T_26; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 564:23 565:14 570:14]
  wire [7:0] _z_result_T_47 = z_result_1 ^ z_result_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 588:32]
  wire [7:0] z_result_4 = z_isResultNaN ? 8'h7f : _z_result_T_47; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 582:23 583:14 588:14]
  wire  z_isResultNaN_5 = _z_isResultNaN_T_4 & _z_isResultNaN_T_9; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 598:34]
  wire [7:0] _GEN_16 = a_data != b_data ? 8'h38 : 8'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 606:42 608:14 610:14]
  wire [7:0] z_result_5 = z_isResultNaN_5 ? 8'h7f : _GEN_16; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 601:23 602:14]
  wire [7:0] _GEN_18 = compareMode == 3'h4 ? z_result_4 : z_result_5; // @[\\src\\main\\scala\\fpu8\\Compare.scala 21:37 22:9 24:9]
  wire [7:0] _GEN_19 = compareMode == 3'h3 ? z_result_3 : _GEN_18; // @[\\src\\main\\scala\\fpu8\\Compare.scala 19:37 20:9]
  wire [7:0] _GEN_20 = compareMode == 3'h2 ? z_result_2 : _GEN_19; // @[\\src\\main\\scala\\fpu8\\Compare.scala 17:37 18:9]
  wire [7:0] _GEN_21 = compareMode == 3'h1 ? z_result_1 : _GEN_20; // @[\\src\\main\\scala\\fpu8\\Compare.scala 15:37 16:9]
  wire [7:0] _GEN_22 = compareMode == 3'h0 ? z_result : _GEN_21; // @[\\src\\main\\scala\\fpu8\\Compare.scala 13:31 14:9]
  assign z = enable ? _GEN_22 : 8'h0; // @[\\src\\main\\scala\\fpu8\\Compare.scala 12:23 27:6]
endmodule
module Convert(
  input        enable, // @[\\src\\main\\scala\\fpu8\\Convert.scala 6:18]
  input  [7:0] a_data, // @[\\src\\main\\scala\\fpu8\\Convert.scala 7:13]
  output [7:0] z // @[\\src\\main\\scala\\fpu8\\Convert.scala 10:13]
);
  wire  _z_fraction_T_1 = a_data[6:3] == 4'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 33:39]
  wire  _z_fraction_T_2 = ~_z_fraction_T_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 617:24]
  wire [3:0] z_fraction = {_z_fraction_T_2,a_data[2:0]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 617:23]
  wire [3:0] _z_leadingZeros_T_8 = {z_fraction[0],z_fraction[1],z_fraction[2],z_fraction[3]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 58:44]
  wire [1:0] _z_leadingZeros_T_13 = _z_leadingZeros_T_8[2] ? 2'h2 : 2'h3; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [1:0] _z_leadingZeros_T_14 = _z_leadingZeros_T_8[1] ? 2'h1 : _z_leadingZeros_T_13; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [1:0] z_shift = _z_leadingZeros_T_8[0] ? 2'h0 : _z_leadingZeros_T_14; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _z_shiftedValue_T_3 = {z_fraction, 1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 63:23]
  wire [5:0] _z_shiftedValue_T_5 = {z_fraction, 2'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 63:23]
  wire [6:0] _z_shiftedValue_T_7 = {z_fraction, 3'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 63:23]
  wire [3:0] _z_shiftedValue_T_10 = 2'h1 == z_shift ? _z_shiftedValue_T_3[3:0] : z_fraction; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [3:0] _z_shiftedValue_T_12 = 2'h2 == z_shift ? _z_shiftedValue_T_5[3:0] : _z_shiftedValue_T_10; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [3:0] z_shiftedFraction = 2'h3 == z_shift ? _z_shiftedValue_T_7[3:0] : _z_shiftedValue_T_12; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [3:0] _GEN_4 = {{2'd0}, z_shift}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 620:40]
  wire [4:0] _z_tempExponent_T_2 = 4'h9 - _GEN_4; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 620:40]
  wire [4:0] _z_tempExponent_T_5 = 4'h8 + a_data[6:3]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 620:54]
  wire [4:0] z_tempExponent = _z_fraction_T_1 ? _z_tempExponent_T_2 : _z_tempExponent_T_5; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 620:27]
  wire [2:0] z_tempFraction = z_shiftedFraction[3:1]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 621:39]
  wire  z_addOne = |a_data[6:3] & &z_shiftedFraction[1:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 623:38]
  wire [2:0] _GEN_5 = {{2'd0}, z_addOne}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 625:40]
  wire [3:0] z_roundedFraction = z_tempFraction + _GEN_5; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 625:40]
  wire [4:0] _z_finalExponent_T_3 = z_tempExponent + 5'h1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 627:83]
  wire [4:0] z_finalExponent = z_roundedFraction[3] ? _z_finalExponent_T_3 : z_tempExponent; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 627:28]
  wire [2:0] z_finalFraction = z_roundedFraction[3] ? z_roundedFraction[3:1] : z_roundedFraction[2:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 628:28]
  wire  _z_T_3 = a_data[2:0] == 3'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 37:44]
  wire  _z_T_4 = _z_fraction_T_1 & _z_T_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 51:26]
  wire  _z_T_7 = a_data[6:3] == 4'hf; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 35:41]
  wire  _z_T_9 = a_data[2:0] == 3'h7; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 39:46]
  wire  _z_T_10 = _z_T_7 & _z_T_9; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 41:30]
  wire  _z_T_11 = ~_z_T_10; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 634:18]
  wire [7:0] _z_result_T_2 = {a_data[7],z_finalExponent,z_finalFraction[1:0]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 635:20]
  wire [7:0] _z_result_T_4 = {a_data[7],5'h0,2'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 637:20]
  wire [7:0] _GEN_0 = _z_T_10 ? 8'h7f : 8'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 638:23 639:14 641:14]
  wire [7:0] _GEN_1 = _z_T_4 & _z_T_11 ? _z_result_T_4 : _GEN_0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 636:31 637:14]
  wire [7:0] z_result = ~_z_T_4 & ~_z_T_10 ? _z_result_T_2 : _GEN_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 634:26 635:14]
  assign z = enable ? z_result : 8'h0; // @[\\src\\main\\scala\\fpu8\\Convert.scala 12:23 13:7 18:7]
endmodule
module GenerateFinalResult(
  input        enable, // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 12:18]
  input        sign, // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 13:16]
  input  [3:0] exponent, // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 14:20]
  input  [2:0] mantissa, // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 15:20]
  input  [1:0] roundingMode, // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 16:24]
  input        overflow, // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 17:20]
  input        saturationMode, // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 18:26]
  input        is0, // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 20:15]
  input        isNaN, // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 21:17]
  output [7:0] z // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 23:13]
);
  wire  _result_T_4 = ~isNaN; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 40:18]
  wire  _result_T_6 = roundingMode == 2'h0; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 42:28]
  wire  _result_T_7 = ~saturationMode; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 42:54]
  wire  _result_T_9 = roundingMode == 2'h1; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 43:26]
  wire  _result_T_10 = roundingMode == 2'h2; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 43:50]
  wire  _result_T_14 = ~sign; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 43:93]
  wire  _result_T_15 = (roundingMode == 2'h1 | roundingMode == 2'h2) & _result_T_7 & ~sign; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 43:85]
  wire  _result_T_16 = roundingMode == 2'h0 & ~saturationMode | _result_T_15; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 42:63]
  wire [7:0] _result_z_T_1 = {sign,4'hf,3'h6}; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 46:19]
  wire [7:0] _GEN_0 = _result_T_9 & sign | _result_T_10 & saturationMode & _result_T_14 ? 8'h7e : 8'h0; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 49:128 50:13 52:13]
  wire [7:0] _GEN_1 = _result_T_9 & saturationMode & _result_T_14 | _result_T_10 & sign ? 8'hfe : _GEN_0; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 47:128 48:13]
  wire [7:0] _GEN_2 = _result_T_6 & saturationMode | roundingMode == 2'h3 & _result_T_7 ? _result_z_T_1 : _GEN_1; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 45:122 46:13]
  wire [7:0] _GEN_3 = _result_T_16 ? 8'h7f : _GEN_2; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 43:103 44:13]
  wire [7:0] _result_z_T_4 = {sign,exponent,mantissa}; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 55:17]
  wire [7:0] _GEN_4 = overflow ? _GEN_3 : _result_z_T_4; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 41:22 55:11]
  wire [7:0] _GEN_5 = isNaN ? 8'h7f : 8'h0; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 59:23 60:9 62:9]
  wire [7:0] _GEN_6 = is0 & _result_T_4 ? 8'h0 : _GEN_5; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 57:31 58:9]
  wire [7:0] result = ~is0 & ~isNaN ? _GEN_4 : _GEN_6; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 40:26]
  assign z = enable ? result : 8'h0; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 31:23 32:7 34:7]
endmodule
module FPU8Generator(
  input        clock,
  input        reset,
  input        enable, // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 9:18]
  input  [7:0] a_data, // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 10:13]
  input  [7:0] b_data, // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 11:13]
  input  [3:0] opCode, // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 12:18]
  input  [1:0] roundingMode, // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 13:24]
  input        saturationMode, // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 14:26]
  output [7:0] z // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 15:13]
);
  wire  addSub_enable; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 17:22]
  wire [7:0] addSub_a_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 17:22]
  wire [7:0] addSub_b_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 17:22]
  wire  addSub_subtract; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 17:22]
  wire [1:0] addSub_roundingMode; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 17:22]
  wire  addSub_sign; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 17:22]
  wire [4:0] addSub_exponent; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 17:22]
  wire [3:0] addSub_fraction; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 17:22]
  wire  addSub_overflow; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 17:22]
  wire  addSub_is0; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 17:22]
  wire  addSub_isNaN; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 17:22]
  wire  multiply_enable; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 19:24]
  wire [7:0] multiply_a_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 19:24]
  wire [7:0] multiply_b_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 19:24]
  wire [1:0] multiply_roundingMode; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 19:24]
  wire  multiply_sign; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 19:24]
  wire [4:0] multiply_exponent; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 19:24]
  wire [3:0] multiply_fraction; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 19:24]
  wire  multiply_overflow; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 19:24]
  wire  multiply_is0; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 19:24]
  wire  multiply_isNaN; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 19:24]
  wire  divide_enable; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 21:22]
  wire [7:0] divide_a_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 21:22]
  wire [7:0] divide_b_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 21:22]
  wire [1:0] divide_roundingMode; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 21:22]
  wire  divide_sign; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 21:22]
  wire [4:0] divide_exponent; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 21:22]
  wire [3:0] divide_fraction; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 21:22]
  wire  divide_overflow; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 21:22]
  wire  divide_is0; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 21:22]
  wire  divide_isNaN; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 21:22]
  wire  compare_enable; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 23:23]
  wire [2:0] compare_compareMode; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 23:23]
  wire [7:0] compare_a_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 23:23]
  wire [7:0] compare_b_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 23:23]
  wire [7:0] compare_z; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 23:23]
  wire  convert_enable; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 25:23]
  wire [7:0] convert_a_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 25:23]
  wire [7:0] convert_z; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 25:23]
  wire  generateFinalResult_enable; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 27:35]
  wire  generateFinalResult_sign; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 27:35]
  wire [3:0] generateFinalResult_exponent; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 27:35]
  wire [2:0] generateFinalResult_mantissa; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 27:35]
  wire [1:0] generateFinalResult_roundingMode; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 27:35]
  wire  generateFinalResult_overflow; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 27:35]
  wire  generateFinalResult_saturationMode; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 27:35]
  wire  generateFinalResult_is0; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 27:35]
  wire  generateFinalResult_isNaN; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 27:35]
  wire [7:0] generateFinalResult_z; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 27:35]
  wire  _addSub_enable_T_2 = opCode == 4'h0 | opCode == 4'h1; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 29:39]
  wire  _multiply_enable_T = opCode == 4'h2; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 35:33]
  wire  _divide_enable_T = opCode == 4'h3; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 40:31]
  wire  _compare_enable_T = opCode == 4'h4; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 45:32]
  wire  _compare_enable_T_1 = opCode == 4'h5; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 45:50]
  wire  _compare_enable_T_3 = opCode == 4'h6; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 45:68]
  wire  _compare_enable_T_5 = opCode == 4'h7; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 45:86]
  wire  _compare_enable_T_7 = opCode == 4'h8; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 45:104]
  wire  _compare_enable_T_10 = opCode == 4'h4 | opCode == 4'h5 | opCode == 4'h6 | opCode == 4'h7 | opCode == 4'h8 |
    opCode == 4'h9; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 45:112]
  wire [2:0] _compare_compareMode_T_5 = _compare_enable_T_7 ? 3'h4 : 3'h5; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 51:14]
  wire [2:0] _compare_compareMode_T_6 = _compare_enable_T_5 ? 3'h3 : _compare_compareMode_T_5; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 50:12]
  wire [2:0] _compare_compareMode_T_7 = _compare_enable_T_3 ? 3'h2 : _compare_compareMode_T_6; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 49:10]
  wire [2:0] _compare_compareMode_T_8 = _compare_enable_T_1 ? 3'h1 : _compare_compareMode_T_7; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 48:8]
  wire  _convert_enable_T = opCode == 4'ha; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 55:32]
  wire [7:0] _GEN_1 = _convert_enable_T ? convert_z : 8'h0; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 114:30 126:7 139:7]
  wire [7:0] _GEN_3 = _compare_enable_T_10 ? compare_z : _GEN_1; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 101:119 113:7]
  wire  _GEN_4 = _divide_enable_T & divide_sign; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 88:30 89:30]
  wire [3:0] _GEN_5 = _divide_enable_T ? divide_exponent[3:0] : 4'h0; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 88:30 90:34]
  wire [2:0] _GEN_6 = _divide_enable_T ? divide_fraction[2:0] : 3'h0; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 88:30 91:34]
  wire [1:0] _GEN_7 = _divide_enable_T ? roundingMode : 2'h0; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 88:30 92:38]
  wire  _GEN_8 = _divide_enable_T & divide_overflow; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 88:30 93:34]
  wire  _GEN_9 = _divide_enable_T & saturationMode; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 88:30 94:40]
  wire  _GEN_11 = _divide_enable_T & divide_is0; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 88:30 96:29]
  wire  _GEN_12 = _divide_enable_T & divide_isNaN; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 88:30 97:31]
  wire [7:0] _GEN_14 = _divide_enable_T ? generateFinalResult_z : _GEN_3; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 88:30 100:7]
  wire  _GEN_15 = _multiply_enable_T ? multiply_sign : _GEN_4; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 75:30 76:30]
  wire [3:0] _GEN_16 = _multiply_enable_T ? multiply_exponent[3:0] : _GEN_5; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 75:30 77:34]
  wire [2:0] _GEN_17 = _multiply_enable_T ? multiply_fraction[2:0] : _GEN_6; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 75:30 78:34]
  wire [1:0] _GEN_18 = _multiply_enable_T ? roundingMode : _GEN_7; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 75:30 79:38]
  wire  _GEN_19 = _multiply_enable_T ? multiply_overflow : _GEN_8; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 75:30 80:34]
  wire  _GEN_20 = _multiply_enable_T ? saturationMode : _GEN_9; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 75:30 81:40]
  wire  _GEN_22 = _multiply_enable_T ? multiply_is0 : _GEN_11; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 75:30 83:29]
  wire  _GEN_23 = _multiply_enable_T ? multiply_isNaN : _GEN_12; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 75:30 84:31]
  wire [7:0] _GEN_25 = _multiply_enable_T ? generateFinalResult_z : _GEN_14; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 75:30 87:7]
  Add addSub ( // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 17:22]
    .enable(addSub_enable),
    .a_data(addSub_a_data),
    .b_data(addSub_b_data),
    .subtract(addSub_subtract),
    .roundingMode(addSub_roundingMode),
    .sign(addSub_sign),
    .exponent(addSub_exponent),
    .fraction(addSub_fraction),
    .overflow(addSub_overflow),
    .is0(addSub_is0),
    .isNaN(addSub_isNaN)
  );
  Multiply multiply ( // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 19:24]
    .enable(multiply_enable),
    .a_data(multiply_a_data),
    .b_data(multiply_b_data),
    .roundingMode(multiply_roundingMode),
    .sign(multiply_sign),
    .exponent(multiply_exponent),
    .fraction(multiply_fraction),
    .overflow(multiply_overflow),
    .is0(multiply_is0),
    .isNaN(multiply_isNaN)
  );
  Divide divide ( // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 21:22]
    .enable(divide_enable),
    .a_data(divide_a_data),
    .b_data(divide_b_data),
    .roundingMode(divide_roundingMode),
    .sign(divide_sign),
    .exponent(divide_exponent),
    .fraction(divide_fraction),
    .overflow(divide_overflow),
    .is0(divide_is0),
    .isNaN(divide_isNaN)
  );
  Compare compare ( // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 23:23]
    .enable(compare_enable),
    .compareMode(compare_compareMode),
    .a_data(compare_a_data),
    .b_data(compare_b_data),
    .z(compare_z)
  );
  Convert convert ( // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 25:23]
    .enable(convert_enable),
    .a_data(convert_a_data),
    .z(convert_z)
  );
  GenerateFinalResult generateFinalResult ( // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 27:35]
    .enable(generateFinalResult_enable),
    .sign(generateFinalResult_sign),
    .exponent(generateFinalResult_exponent),
    .mantissa(generateFinalResult_mantissa),
    .roundingMode(generateFinalResult_roundingMode),
    .overflow(generateFinalResult_overflow),
    .saturationMode(generateFinalResult_saturationMode),
    .is0(generateFinalResult_is0),
    .isNaN(generateFinalResult_isNaN),
    .z(generateFinalResult_z)
  );
  assign z = _addSub_enable_T_2 ? generateFinalResult_z : _GEN_25; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 62:42 74:7]
  assign addSub_enable = (opCode == 4'h0 | opCode == 4'h1) & enable; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 29:23]
  assign addSub_a_data = a_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 30:12]
  assign addSub_b_data = b_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 31:12]
  assign addSub_subtract = opCode == 4'h1; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 32:33]
  assign addSub_roundingMode = roundingMode; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 33:23]
  assign multiply_enable = opCode == 4'h2 & enable; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 35:25]
  assign multiply_a_data = a_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 36:14]
  assign multiply_b_data = b_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 37:14]
  assign multiply_roundingMode = roundingMode; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 38:25]
  assign divide_enable = opCode == 4'h3 & enable; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 40:23]
  assign divide_a_data = a_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 41:12]
  assign divide_b_data = b_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 42:12]
  assign divide_roundingMode = roundingMode; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 43:23]
  assign compare_enable = (opCode == 4'h4 | opCode == 4'h5 | opCode == 4'h6 | opCode == 4'h7 | opCode == 4'h8 | opCode
     == 4'h9) & enable; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 45:24]
  assign compare_compareMode = _compare_enable_T ? 3'h0 : _compare_compareMode_T_8; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 47:29]
  assign compare_a_data = a_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 52:13]
  assign compare_b_data = b_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 53:13]
  assign convert_enable = opCode == 4'ha & enable; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 55:24]
  assign convert_a_data = a_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 56:13]
  assign generateFinalResult_enable = enable; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 60:30]
  assign generateFinalResult_sign = _addSub_enable_T_2 ? addSub_sign : _GEN_15; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 62:42 63:30]
  assign generateFinalResult_exponent = _addSub_enable_T_2 ? addSub_exponent[3:0] : _GEN_16; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 62:42 64:34]
  assign generateFinalResult_mantissa = _addSub_enable_T_2 ? addSub_fraction[2:0] : _GEN_17; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 62:42 65:34]
  assign generateFinalResult_roundingMode = _addSub_enable_T_2 ? roundingMode : _GEN_18; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 62:42 66:38]
  assign generateFinalResult_overflow = _addSub_enable_T_2 ? addSub_overflow : _GEN_19; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 62:42 67:34]
  assign generateFinalResult_saturationMode = _addSub_enable_T_2 ? saturationMode : _GEN_20; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 62:42 68:40]
  assign generateFinalResult_is0 = _addSub_enable_T_2 ? addSub_is0 : _GEN_22; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 62:42 70:29]
  assign generateFinalResult_isNaN = _addSub_enable_T_2 ? addSub_isNaN : _GEN_23; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 62:42 71:31]
endmodule
