module Add(
  input        enable, // @[\\src\\main\\scala\\fpu8\\Add.scala 10:18]
  input  [7:0] a_data, // @[\\src\\main\\scala\\fpu8\\Add.scala 11:13]
  input  [7:0] b_data, // @[\\src\\main\\scala\\fpu8\\Add.scala 12:13]
  input        subtract, // @[\\src\\main\\scala\\fpu8\\Add.scala 13:20]
  input  [1:0] roundingMode, // @[\\src\\main\\scala\\fpu8\\Add.scala 14:24]
  output       sign, // @[\\src\\main\\scala\\fpu8\\Add.scala 15:16]
  output [4:0] exponent, // @[\\src\\main\\scala\\fpu8\\Add.scala 16:20]
  output [3:0] fraction, // @[\\src\\main\\scala\\fpu8\\Add.scala 17:20]
  output [4:0] status // @[\\src\\main\\scala\\fpu8\\Add.scala 19:18]
);
  wire  compare = a_data[6:0] > b_data[6:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 29:77]
  wire [7:0] greaterOperand_data = compare ? a_data : b_data; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 131:29]
  wire [7:0] smallerOperand_data = compare ? b_data : a_data; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 132:29]
  wire  resultSign = compare ? a_data[7] : b_data[7] ^ subtract; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 133:19]
  wire  subtraction = subtract ^ greaterOperand_data[7] ^ smallerOperand_data[7]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 134:54]
  wire [3:0] exponent_1 = greaterOperand_data[6:3]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 25:28]
  wire  _greaterOperandFraction_T_1 = exponent_1 == 4'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 35:39]
  wire  _greaterOperandFraction_T_2 = ~_greaterOperandFraction_T_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 136:38]
  wire  _smallerOperandFraction_T_1 = smallerOperand_data[6:3] == 4'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 35:39]
  wire  _smallerOperandFraction_T_2 = ~_smallerOperandFraction_T_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 137:38]
  wire  isOnlySmallerDenormalized = _greaterOperandFraction_T_2 & _smallerOperandFraction_T_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 138:60]
  wire [3:0] _shift_T_2 = exponent_1 - 4'h1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 141:31]
  wire [3:0] _shift_T_6 = exponent_1 - smallerOperand_data[6:3]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 142:31]
  wire [3:0] shift = isOnlySmallerDenormalized ? _shift_T_2 : _shift_T_6; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 139:20]
  wire  _shiftedFraction_shifted_T = shift >= 4'h6; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 147:15]
  wire [9:0] _shiftedFraction_shifted_T_1 = {6'h0,_smallerOperandFraction_T_2,smallerOperand_data[2:0]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 148:12]
  wire [9:0] _shiftedFraction_shifted_T_2 = {_smallerOperandFraction_T_2,smallerOperand_data[2:0],6'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 149:12]
  wire [9:0] _shiftedFraction_shifted_T_3 = _shiftedFraction_shifted_T_2 >> shift; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 149:54]
  wire [9:0] shiftedFraction_shifted = _shiftedFraction_shifted_T ? _shiftedFraction_shifted_T_1 :
    _shiftedFraction_shifted_T_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 146:24]
  wire [6:0] smallerOperandFraction_1 = {shiftedFraction_shifted[9:4],|shiftedFraction_shifted[3:0]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 151:10]
  wire [6:0] greaterOperandFraction_1 = {_greaterOperandFraction_T_2,greaterOperand_data[2:0],3'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 153:45]
  wire  _isResultNaN_T_1 = a_data[6:3] == 4'hf; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 37:41]
  wire  _isResultNaN_T_3 = a_data[2:0] == 3'h7; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 41:46]
  wire  _isResultNaN_T_4 = _isResultNaN_T_1 & _isResultNaN_T_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 43:30]
  wire  _isResultNaN_T_6 = b_data[6:3] == 4'hf; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 37:41]
  wire  _isResultNaN_T_8 = b_data[2:0] == 3'h7; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 41:46]
  wire  _isResultNaN_T_9 = _isResultNaN_T_6 & _isResultNaN_T_8; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 43:30]
  wire  isResultNaN = _isResultNaN_T_4 | _isResultNaN_T_9; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 416:37]
  wire  _isResult0_T_2 = a_data[6:0] == b_data[6:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 33:77]
  wire  isResult0 = _isResult0_T_2 & subtraction & ~isResultNaN; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 424:85]
  wire [7:0] _calculatedValue_T_1 = greaterOperandFraction_1 - smallerOperandFraction_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 429:32]
  wire [7:0] _calculatedValue_T_3 = greaterOperandFraction_1 + smallerOperandFraction_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 430:32]
  wire [7:0] calculatedValue = subtraction ? _calculatedValue_T_1 : _calculatedValue_T_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 428:32]
  wire [6:0] _leadingZeros_T_17 = {calculatedValue[0],calculatedValue[1],calculatedValue[2],calculatedValue[3],
    calculatedValue[4],calculatedValue[5],calculatedValue[6]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 60:44]
  wire [2:0] _leadingZeros_T_25 = _leadingZeros_T_17[5] ? 3'h5 : 3'h6; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] _leadingZeros_T_26 = _leadingZeros_T_17[4] ? 3'h4 : _leadingZeros_T_25; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] _leadingZeros_T_27 = _leadingZeros_T_17[3] ? 3'h3 : _leadingZeros_T_26; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] _leadingZeros_T_28 = _leadingZeros_T_17[2] ? 3'h2 : _leadingZeros_T_27; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] _leadingZeros_T_29 = _leadingZeros_T_17[1] ? 3'h1 : _leadingZeros_T_28; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] shift_1 = _leadingZeros_T_17[0] ? 3'h0 : _leadingZeros_T_29; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [7:0] _shiftedValue_T_3 = {calculatedValue[6:0], 1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 65:23]
  wire [8:0] _shiftedValue_T_5 = {calculatedValue[6:0], 2'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 65:23]
  wire [9:0] _shiftedValue_T_7 = {calculatedValue[6:0], 3'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 65:23]
  wire [10:0] _shiftedValue_T_9 = {calculatedValue[6:0], 4'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 65:23]
  wire [11:0] _shiftedValue_T_11 = {calculatedValue[6:0], 5'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 65:23]
  wire [12:0] _shiftedValue_T_13 = {calculatedValue[6:0], 6'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 65:23]
  wire [6:0] _shiftedValue_T_18 = 3'h1 == shift_1 ? _shiftedValue_T_3[6:0] : calculatedValue[6:0]; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [6:0] _shiftedValue_T_20 = 3'h2 == shift_1 ? _shiftedValue_T_5[6:0] : _shiftedValue_T_18; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [6:0] _shiftedValue_T_22 = 3'h3 == shift_1 ? _shiftedValue_T_7[6:0] : _shiftedValue_T_20; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [6:0] _shiftedValue_T_24 = 3'h4 == shift_1 ? _shiftedValue_T_9[6:0] : _shiftedValue_T_22; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [6:0] _shiftedValue_T_26 = 3'h5 == shift_1 ? _shiftedValue_T_11[6:0] : _shiftedValue_T_24; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [6:0] shiftedCalcValue = 3'h6 == shift_1 ? _shiftedValue_T_13[6:0] : _shiftedValue_T_26; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _T_1 = &exponent_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 277:19]
  wire [3:0] _tempExponent_T_1 = exponent_1 + 4'h1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 281:32]
  wire [6:0] _tempFraction_T_3 = {calculatedValue[7:2],|calculatedValue[1:0]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 282:26]
  wire [3:0] _GEN_12 = {{1'd0}, shift_1}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 283:25]
  wire [3:0] _tempExponent_T_3 = exponent_1 - _GEN_12; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 284:32]
  wire [21:0] _GEN_5 = {{15'd0}, calculatedValue[6:0]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 289:47]
  wire [21:0] _tempFraction_T_7 = _GEN_5 << _shift_T_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 289:47]
  wire [21:0] _GEN_0 = exponent_1 > 4'h0 ? _tempFraction_T_7 : {{15'd0}, calculatedValue[6:0]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 288:28 289:22 291:22]
  wire [3:0] _GEN_1 = exponent_1 > _GEN_12 & shiftedCalcValue[6] ? _tempExponent_T_3 : 4'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 283:57 284:20 287:20]
  wire [21:0] _GEN_2 = exponent_1 > _GEN_12 & shiftedCalcValue[6] ? {{15'd0}, shiftedCalcValue} : _GEN_0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 283:57 285:20]
  wire [3:0] _GEN_3 = ~_T_1 & calculatedValue[7] ? _tempExponent_T_1 : _GEN_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 280:54 281:20]
  wire [21:0] _GEN_4 = ~_T_1 & calculatedValue[7] ? {{15'd0}, _tempFraction_T_3} : _GEN_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 280:54 282:20]
  wire [3:0] tempExponent = &exponent_1 & calculatedValue[7] ? exponent_1 : _GEN_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 277:47 278:20]
  wire [21:0] _GEN_6 = &exponent_1 & calculatedValue[7] ? 22'h7f : _GEN_4; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 277:47 279:20]
  wire [6:0] tempFraction = _GEN_6[6:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 275:28]
  wire  _addOne_T_2 = roundingMode == 2'h0 & tempFraction[2]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 236:42]
  wire  _addOne_T_17 = _addOne_T_2 & ~tempFraction[1] & ~tempFraction[0] & tempFraction[3]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 237:90]
  wire  _addOne_T_18 = roundingMode == 2'h0 & tempFraction[2] & (tempFraction[1] | tempFraction[0]) | _addOne_T_17; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 236:102]
  wire  _addOne_T_24 = tempFraction[2] | tempFraction[1] | tempFraction[0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 238:70]
  wire  _addOne_T_27 = roundingMode == 2'h1 & (tempFraction[2] | tempFraction[1] | tempFraction[0]) & resultSign; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 238:90]
  wire  _addOne_T_28 = _addOne_T_18 | _addOne_T_27; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 237:110]
  wire  _addOne_T_38 = roundingMode == 2'h2 & _addOne_T_24 & ~resultSign; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 239:90]
  wire  addOne = _addOne_T_28 | _addOne_T_38; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 238:106]
  wire [3:0] _GEN_14 = {{3'd0}, addOne}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 241:66]
  wire [4:0] roundedFraction = tempFraction[6:3] + _GEN_14; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 241:66]
  wire [3:0] resultFraction = roundedFraction[4] ? roundedFraction[4:1] : roundedFraction[3:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 243:28]
  wire [3:0] _finalExponent_T_7 = tempExponent + 4'h1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 247:20]
  wire [3:0] resultExponent = roundedFraction[4] | roundedFraction[3] & tempExponent == 4'h0 ? _finalExponent_T_7 :
    tempExponent; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 246:28]
  wire  _overflow_T_9 = tempExponent >= 4'hf & tempFraction[6:3] == 4'hf; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 252:42]
  wire  overflow = resultExponent == 4'hf & resultFraction == 4'hf | _overflow_T_9; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 251:134]
  wire [4:0] resultStatus = {overflow,resultExponent == 4'h0,isResultNaN,1'h0,isResult0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 434:23]
  wire [3:0] _GEN_8 = enable ? resultExponent : 4'h0; // @[\\src\\main\\scala\\fpu8\\Add.scala 24:24 26:14 32:14]
  assign sign = enable & resultSign; // @[\\src\\main\\scala\\fpu8\\Add.scala 24:24 25:10 31:10]
  assign exponent = {{1'd0}, _GEN_8};
  assign fraction = enable ? resultFraction : 4'h0; // @[\\src\\main\\scala\\fpu8\\Add.scala 24:24 27:14 33:14]
  assign status = enable ? resultStatus : 5'h0; // @[\\src\\main\\scala\\fpu8\\Add.scala 24:24 28:12 34:12]
endmodule
module Multiply(
  input        enable, // @[\\src\\main\\scala\\fpu8\\Multiply.scala 10:18]
  input  [7:0] a_data, // @[\\src\\main\\scala\\fpu8\\Multiply.scala 11:13]
  input  [7:0] b_data, // @[\\src\\main\\scala\\fpu8\\Multiply.scala 12:13]
  input  [1:0] roundingMode, // @[\\src\\main\\scala\\fpu8\\Multiply.scala 13:24]
  output       sign, // @[\\src\\main\\scala\\fpu8\\Multiply.scala 14:16]
  output [4:0] exponent, // @[\\src\\main\\scala\\fpu8\\Multiply.scala 15:20]
  output [3:0] fraction, // @[\\src\\main\\scala\\fpu8\\Multiply.scala 16:20]
  output [4:0] status // @[\\src\\main\\scala\\fpu8\\Multiply.scala 18:18]
);
  wire  _isResultNaN_T_1 = a_data[6:3] == 4'hf; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 37:41]
  wire  _isResultNaN_T_3 = a_data[2:0] == 3'h7; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 41:46]
  wire  _isResultNaN_T_4 = _isResultNaN_T_1 & _isResultNaN_T_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 43:30]
  wire  _isResultNaN_T_6 = b_data[6:3] == 4'hf; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 37:41]
  wire  _isResultNaN_T_8 = b_data[2:0] == 3'h7; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 41:46]
  wire  _isResultNaN_T_9 = _isResultNaN_T_6 & _isResultNaN_T_8; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 43:30]
  wire  isResultNaN = _isResultNaN_T_4 | _isResultNaN_T_9; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 446:37]
  wire  _isResult0_T_1 = a_data[6:3] == 4'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 35:39]
  wire  _isResult0_T_3 = a_data[2:0] == 3'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 39:44]
  wire  _isResult0_T_4 = _isResult0_T_1 & _isResult0_T_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 53:26]
  wire  _isResult0_T_15 = b_data[6:3] == 4'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 35:39]
  wire  _isResult0_T_17 = b_data[2:0] == 3'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 39:44]
  wire  _isResult0_T_18 = _isResult0_T_15 & _isResult0_T_17; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 53:26]
  wire  isResult0 = _isResult0_T_4 & ~_isResultNaN_T_9 | _isResult0_T_18 & ~_isResultNaN_T_4; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 454:80]
  wire  resultSign = a_data[7] ^ b_data[7]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 158:26]
  wire [5:0] _exponent_T_11 = {2'h0,a_data[6:3]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 164:16]
  wire [5:0] _exponent_T_13 = {2'h0,b_data[6:3]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 164:47]
  wire [5:0] _exponent_T_15 = _exponent_T_11 + _exponent_T_13; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 164:42]
  wire [5:0] _exponent_T_17 = _exponent_T_15 - 6'h6; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 164:74]
  wire [5:0] _exponent_T_25 = _exponent_T_15 - 6'h7; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 165:74]
  wire [5:0] _exponent_T_26 = _isResult0_T_1 ^ _isResult0_T_15 ? _exponent_T_17 : _exponent_T_25; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 163:14]
  wire [5:0] exponent_1 = _isResult0_T_1 & _isResult0_T_15 ? 6'h34 : _exponent_T_26; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 161:12]
  wire  _firstOperandFraction_T_2 = ~_isResult0_T_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 173:36]
  wire [3:0] firstOperandFraction = {_firstOperandFraction_T_2,a_data[2:0]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 173:35]
  wire  _secondOperandFraction_T_2 = ~_isResult0_T_15; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 174:37]
  wire [3:0] secondOperandFraction = {_secondOperandFraction_T_2,b_data[2:0]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 174:36]
  wire [3:0] product_partialProducts_compare = secondOperandFraction[0] ? 4'hf : 4'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 103:24]
  wire [3:0] product_partialProducts_0 = firstOperandFraction & product_partialProducts_compare; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:11]
  wire [3:0] product_partialProducts_compare_1 = secondOperandFraction[1] ? 4'hf : 4'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 103:24]
  wire [3:0] _product_partialProducts_T_1 = firstOperandFraction & product_partialProducts_compare_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:11]
  wire [4:0] product_partialProducts_1 = {_product_partialProducts_T_1, 1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:22]
  wire [3:0] product_partialProducts_compare_2 = secondOperandFraction[2] ? 4'hf : 4'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 103:24]
  wire [3:0] _product_partialProducts_T_2 = firstOperandFraction & product_partialProducts_compare_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:11]
  wire [5:0] product_partialProducts_2 = {_product_partialProducts_T_2, 2'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:22]
  wire [3:0] product_partialProducts_compare_3 = secondOperandFraction[3] ? 4'hf : 4'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 103:24]
  wire [3:0] _product_partialProducts_T_3 = firstOperandFraction & product_partialProducts_compare_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:11]
  wire [6:0] product_partialProducts_3 = {_product_partialProducts_T_3, 3'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:22]
  wire [4:0] _GEN_12 = {{1'd0}, product_partialProducts_0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 114:34]
  wire [5:0] _product_partialSums_T = _GEN_12 + product_partialProducts_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 114:34]
  wire [6:0] product_partialSums_0 = _product_partialSums_T + product_partialProducts_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 114:39]
  wire [7:0] product = product_partialSums_0 + product_partialProducts_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 111:15]
  wire [6:0] _leadingZeros_T_17 = {product[0],product[1],product[2],product[3],product[4],product[5],product[6]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 60:44]
  wire [2:0] _leadingZeros_T_25 = _leadingZeros_T_17[5] ? 3'h5 : 3'h6; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] _leadingZeros_T_26 = _leadingZeros_T_17[4] ? 3'h4 : _leadingZeros_T_25; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] _leadingZeros_T_27 = _leadingZeros_T_17[3] ? 3'h3 : _leadingZeros_T_26; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] _leadingZeros_T_28 = _leadingZeros_T_17[2] ? 3'h2 : _leadingZeros_T_27; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] _leadingZeros_T_29 = _leadingZeros_T_17[1] ? 3'h1 : _leadingZeros_T_28; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] shift = _leadingZeros_T_17[0] ? 3'h0 : _leadingZeros_T_29; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [7:0] _shiftedValue_T_3 = {product[6:0], 1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 65:23]
  wire [8:0] _shiftedValue_T_5 = {product[6:0], 2'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 65:23]
  wire [9:0] _shiftedValue_T_7 = {product[6:0], 3'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 65:23]
  wire [10:0] _shiftedValue_T_9 = {product[6:0], 4'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 65:23]
  wire [11:0] _shiftedValue_T_11 = {product[6:0], 5'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 65:23]
  wire [12:0] _shiftedValue_T_13 = {product[6:0], 6'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 65:23]
  wire [6:0] _shiftedValue_T_18 = 3'h1 == shift ? _shiftedValue_T_3[6:0] : product[6:0]; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [6:0] _shiftedValue_T_20 = 3'h2 == shift ? _shiftedValue_T_5[6:0] : _shiftedValue_T_18; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [6:0] _shiftedValue_T_22 = 3'h3 == shift ? _shiftedValue_T_7[6:0] : _shiftedValue_T_20; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [6:0] _shiftedValue_T_24 = 3'h4 == shift ? _shiftedValue_T_9[6:0] : _shiftedValue_T_22; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [6:0] _shiftedValue_T_26 = 3'h5 == shift ? _shiftedValue_T_11[6:0] : _shiftedValue_T_24; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [6:0] shiftedCalcValue = 3'h6 == shift ? _shiftedValue_T_13[6:0] : _shiftedValue_T_26; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [5:0] exponentShiftRight = 6'h0 - exponent_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 307:55]
  wire [5:0] exponentShiftLeft = exponent_1 - 6'h1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 310:35]
  wire  _T_2 = ~exponent_1[5]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 316:10]
  wire  _T_5 = ~exponent_1[5] & exponent_1[4:0] >= 5'hf; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 316:40]
  wire  _T_12 = _T_2 & exponent_1[4:0] < 5'hf; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 320:46]
  wire [4:0] _tempExponent_T_2 = exponent_1[4:0] + 5'h1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 322:38]
  wire [6:0] _tempFraction_T_3 = {product[7:2],|product[1:0]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 323:26]
  wire [4:0] _GEN_13 = {{2'd0}, shift}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 324:78]
  wire  _T_19 = _T_2 & exponent_1[4:0] > _GEN_13; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 324:46]
  wire [4:0] _tempExponent_T_5 = exponent_1[4:0] - _GEN_13; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 326:51]
  wire [6:0] _tempFraction_T_27 = 6'h0 == exponentShiftLeft ? product[6:0] : product[6:0]; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [6:0] _tempFraction_T_29 = 6'h1 == exponentShiftLeft ? _shiftedValue_T_3[6:0] : _tempFraction_T_27; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [6:0] _tempFraction_T_31 = 6'h2 == exponentShiftLeft ? _shiftedValue_T_5[6:0] : _tempFraction_T_29; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [6:0] _tempFraction_T_33 = 6'h3 == exponentShiftLeft ? _shiftedValue_T_7[6:0] : _tempFraction_T_31; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [6:0] _tempFraction_T_35 = 6'h4 == exponentShiftLeft ? _shiftedValue_T_9[6:0] : _tempFraction_T_33; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [6:0] _tempFraction_T_37 = 6'h5 == exponentShiftLeft ? _shiftedValue_T_11[6:0] : _tempFraction_T_35; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [6:0] _tempFraction_T_39 = 6'h6 == exponentShiftLeft ? _shiftedValue_T_13[6:0] : _tempFraction_T_37; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [6:0] _tempFraction_T_44 = _tempFraction_T_3 >> exponentShiftRight; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 338:110]
  wire [6:0] _GEN_0 = _T_2 & exponent_1[4:0] > 5'h0 ? _tempFraction_T_39 : _tempFraction_T_44; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 330:82 332:22 338:22]
  wire [4:0] _GEN_1 = _T_19 & shiftedCalcValue[6] ? _tempExponent_T_5 : 5'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 325:55 326:20 329:20]
  wire [6:0] _GEN_2 = _T_19 & shiftedCalcValue[6] ? shiftedCalcValue : _GEN_0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 325:55 327:20]
  wire [4:0] _GEN_3 = _T_12 & product[7] ? _tempExponent_T_2 : _GEN_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 321:54 322:20]
  wire [6:0] _GEN_4 = _T_12 & product[7] ? _tempFraction_T_3 : _GEN_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 321:54 323:20]
  wire [4:0] tempExponent = _T_5 & product[7] ? 5'hf : _GEN_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 317:54 318:20]
  wire [6:0] tempFraction = _T_5 & product[7] ? 7'h7f : _GEN_4; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 317:54 319:20]
  wire  _addOne_T_2 = roundingMode == 2'h0 & tempFraction[2]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 236:42]
  wire  _addOne_T_17 = _addOne_T_2 & ~tempFraction[1] & ~tempFraction[0] & tempFraction[3]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 237:90]
  wire  _addOne_T_18 = roundingMode == 2'h0 & tempFraction[2] & (tempFraction[1] | tempFraction[0]) | _addOne_T_17; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 236:102]
  wire  _addOne_T_24 = tempFraction[2] | tempFraction[1] | tempFraction[0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 238:70]
  wire  _addOne_T_27 = roundingMode == 2'h1 & (tempFraction[2] | tempFraction[1] | tempFraction[0]) & resultSign; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 238:90]
  wire  _addOne_T_28 = _addOne_T_18 | _addOne_T_27; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 237:110]
  wire  _addOne_T_38 = roundingMode == 2'h2 & _addOne_T_24 & ~resultSign; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 239:90]
  wire  addOne = _addOne_T_28 | _addOne_T_38; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 238:106]
  wire [3:0] _GEN_15 = {{3'd0}, addOne}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 241:66]
  wire [4:0] roundedFraction = tempFraction[6:3] + _GEN_15; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 241:66]
  wire [3:0] resultFraction = roundedFraction[4] ? roundedFraction[4:1] : roundedFraction[3:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 243:28]
  wire [4:0] _finalExponent_T_7 = tempExponent + 5'h1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 247:20]
  wire [4:0] resultExponent = roundedFraction[4] | roundedFraction[3] & tempExponent == 5'h0 ? _finalExponent_T_7 :
    tempExponent; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 246:28]
  wire  _overflow_T_9 = tempExponent >= 5'hf & tempFraction[6:3] == 4'hf; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 252:42]
  wire  overflow = resultExponent > 5'hf | resultExponent[3:0] == 4'hf & resultFraction == 4'hf | _overflow_T_9; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 251:134]
  wire [4:0] resultStatus = {overflow,resultExponent == 5'h0,isResultNaN,1'h0,isResult0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 464:23]
  assign sign = enable & resultSign; // @[\\src\\main\\scala\\fpu8\\Multiply.scala 23:24 24:10 30:10]
  assign exponent = enable ? resultExponent : 5'h0; // @[\\src\\main\\scala\\fpu8\\Multiply.scala 23:24 25:14 31:14]
  assign fraction = enable ? resultFraction : 4'h0; // @[\\src\\main\\scala\\fpu8\\Multiply.scala 23:24 26:14 32:14]
  assign status = enable ? resultStatus : 5'h0; // @[\\src\\main\\scala\\fpu8\\Multiply.scala 23:24 27:12 33:12]
endmodule
module Divide(
  input        enable, // @[\\src\\main\\scala\\fpu8\\Divide.scala 10:18]
  input  [7:0] a_data, // @[\\src\\main\\scala\\fpu8\\Divide.scala 11:13]
  input  [7:0] b_data, // @[\\src\\main\\scala\\fpu8\\Divide.scala 12:13]
  input  [1:0] roundingMode, // @[\\src\\main\\scala\\fpu8\\Divide.scala 13:24]
  output       sign, // @[\\src\\main\\scala\\fpu8\\Divide.scala 14:16]
  output [4:0] exponent, // @[\\src\\main\\scala\\fpu8\\Divide.scala 15:20]
  output [3:0] fraction, // @[\\src\\main\\scala\\fpu8\\Divide.scala 16:20]
  output [4:0] status // @[\\src\\main\\scala\\fpu8\\Divide.scala 18:18]
);
  wire  _isResultNaN_T_1 = a_data[6:3] == 4'hf; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 37:41]
  wire  _isResultNaN_T_3 = a_data[2:0] == 3'h7; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 41:46]
  wire  _isResultNaN_T_4 = _isResultNaN_T_1 & _isResultNaN_T_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 43:30]
  wire  _isResultNaN_T_6 = b_data[6:3] == 4'hf; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 37:41]
  wire  _isResultNaN_T_8 = b_data[2:0] == 3'h7; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 41:46]
  wire  _isResultNaN_T_9 = _isResultNaN_T_6 & _isResultNaN_T_8; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 43:30]
  wire  _isResultNaN_T_12 = b_data[6:3] == 4'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 35:39]
  wire  _isResultNaN_T_14 = b_data[2:0] == 3'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 39:44]
  wire  _isResultNaN_T_15 = _isResultNaN_T_12 & _isResultNaN_T_14; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 53:26]
  wire  isResultNaN = _isResultNaN_T_4 | _isResultNaN_T_9 | _isResultNaN_T_15; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 476:40]
  wire  _isResult0_T_1 = a_data[6:3] == 4'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 35:39]
  wire  _isResult0_T_3 = a_data[2:0] == 3'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 39:44]
  wire  _isResult0_T_4 = _isResult0_T_1 & _isResult0_T_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 53:26]
  wire  isResult0 = _isResult0_T_4 & ~_isResultNaN_T_15 & ~_isResultNaN_T_9; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 487:37]
  wire  resultSign = a_data[7] ^ b_data[7]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 180:26]
  wire [3:0] _tempDividendFraction_T_3 = {a_data[2:0],1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 182:10]
  wire [3:0] _tempDividendFraction_T_5 = {1'h1,a_data[2:0]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 183:10]
  wire [3:0] tempDividendFraction = _isResult0_T_1 ? _tempDividendFraction_T_3 : _tempDividendFraction_T_5; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 181:35]
  wire [3:0] _tempDivisorFraction_T_3 = {b_data[2:0],1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 186:10]
  wire [3:0] _tempDivisorFraction_T_5 = {1'h1,b_data[2:0]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 187:10]
  wire [3:0] tempDivisorFraction = _isResultNaN_T_12 ? _tempDivisorFraction_T_3 : _tempDivisorFraction_T_5; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 185:34]
  wire [5:0] _tempExponent_T_1 = {2'h0,a_data[6:3]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 189:27]
  wire [5:0] _tempExponent_T_3 = {2'h0,b_data[6:3]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 190:10]
  wire [5:0] _tempExponent_T_5 = _tempExponent_T_1 - _tempExponent_T_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 189:53]
  wire [5:0] tempExponent = _tempExponent_T_5 + 6'h7; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 190:37]
  wire [3:0] _leadingZeros_T_8 = {tempDividendFraction[0],tempDividendFraction[1],tempDividendFraction[2],
    tempDividendFraction[3]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 60:44]
  wire [1:0] _leadingZeros_T_13 = _leadingZeros_T_8[2] ? 2'h2 : 2'h3; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [1:0] _leadingZeros_T_14 = _leadingZeros_T_8[1] ? 2'h1 : _leadingZeros_T_13; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [1:0] dividendShift = _leadingZeros_T_8[0] ? 2'h0 : _leadingZeros_T_14; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _shiftedValue_T_3 = {tempDividendFraction, 1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 65:23]
  wire [5:0] _shiftedValue_T_5 = {tempDividendFraction, 2'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 65:23]
  wire [6:0] _shiftedValue_T_7 = {tempDividendFraction, 3'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 65:23]
  wire [3:0] _shiftedValue_T_10 = 2'h1 == dividendShift ? _shiftedValue_T_3[3:0] : tempDividendFraction; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [3:0] _shiftedValue_T_12 = 2'h2 == dividendShift ? _shiftedValue_T_5[3:0] : _shiftedValue_T_10; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [3:0] dividendFraction = 2'h3 == dividendShift ? _shiftedValue_T_7[3:0] : _shiftedValue_T_12; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [3:0] _leadingZeros_T_24 = {tempDivisorFraction[0],tempDivisorFraction[1],tempDivisorFraction[2],
    tempDivisorFraction[3]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 60:44]
  wire [1:0] _leadingZeros_T_29 = _leadingZeros_T_24[2] ? 2'h2 : 2'h3; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [1:0] _leadingZeros_T_30 = _leadingZeros_T_24[1] ? 2'h1 : _leadingZeros_T_29; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [1:0] divisorShift = _leadingZeros_T_24[0] ? 2'h0 : _leadingZeros_T_30; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _shiftedValue_T_18 = {tempDivisorFraction, 1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 65:23]
  wire [5:0] _shiftedValue_T_20 = {tempDivisorFraction, 2'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 65:23]
  wire [6:0] _shiftedValue_T_22 = {tempDivisorFraction, 3'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 65:23]
  wire [3:0] _shiftedValue_T_25 = 2'h1 == divisorShift ? _shiftedValue_T_18[3:0] : tempDivisorFraction; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [3:0] _shiftedValue_T_27 = 2'h2 == divisorShift ? _shiftedValue_T_20[3:0] : _shiftedValue_T_25; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [3:0] divisorFraction = 2'h3 == divisorShift ? _shiftedValue_T_22[3:0] : _shiftedValue_T_27; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [5:0] _GEN_20 = {{4'd0}, dividendShift}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 197:33]
  wire [5:0] _exponent_T_1 = tempExponent - _GEN_20; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 197:33]
  wire [5:0] _GEN_21 = {{4'd0}, divisorShift}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 197:49]
  wire [5:0] exponent_1 = _exponent_T_1 + _GEN_21; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 197:49]
  wire [3:0] _GEN_1 = 3'h1 == divisorFraction[2:0] ? 4'hc : 4'he; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 205:{24,24}]
  wire [3:0] _GEN_2 = 3'h2 == divisorFraction[2:0] ? 4'ha : _GEN_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 205:{24,24}]
  wire [3:0] _GEN_3 = 3'h3 == divisorFraction[2:0] ? 4'h8 : _GEN_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 205:{24,24}]
  wire [3:0] _GEN_4 = 3'h4 == divisorFraction[2:0] ? 4'h6 : _GEN_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 205:{24,24}]
  wire [3:0] _GEN_5 = 3'h5 == divisorFraction[2:0] ? 4'h4 : _GEN_4; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 205:{24,24}]
  wire [3:0] _GEN_6 = 3'h6 == divisorFraction[2:0] ? 4'h2 : _GEN_5; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 205:{24,24}]
  wire [3:0] _GEN_7 = 3'h7 == divisorFraction[2:0] ? 4'h0 : _GEN_6; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 205:{24,24}]
  wire [5:0] quotient_initGuess = {2'h1,_GEN_7}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 205:24]
  wire [5:0] quotient_secondGuess_firstStep_partialProducts_compare = divisorFraction[0] ? 6'h3f : 6'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 103:24]
  wire [5:0] quotient_secondGuess_firstStep_partialProducts_0 = quotient_initGuess &
    quotient_secondGuess_firstStep_partialProducts_compare; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:11]
  wire [5:0] quotient_secondGuess_firstStep_partialProducts_compare_1 = divisorFraction[1] ? 6'h3f : 6'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 103:24]
  wire [5:0] _quotient_secondGuess_firstStep_partialProducts_T_1 = quotient_initGuess &
    quotient_secondGuess_firstStep_partialProducts_compare_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:11]
  wire [6:0] quotient_secondGuess_firstStep_partialProducts_1 = {_quotient_secondGuess_firstStep_partialProducts_T_1
    , 1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:22]
  wire [5:0] quotient_secondGuess_firstStep_partialProducts_compare_2 = divisorFraction[2] ? 6'h3f : 6'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 103:24]
  wire [5:0] _quotient_secondGuess_firstStep_partialProducts_T_2 = quotient_initGuess &
    quotient_secondGuess_firstStep_partialProducts_compare_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:11]
  wire [7:0] quotient_secondGuess_firstStep_partialProducts_2 = {_quotient_secondGuess_firstStep_partialProducts_T_2
    , 2'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:22]
  wire [5:0] quotient_secondGuess_firstStep_partialProducts_compare_3 = divisorFraction[3] ? 6'h3f : 6'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 103:24]
  wire [5:0] _quotient_secondGuess_firstStep_partialProducts_T_3 = quotient_initGuess &
    quotient_secondGuess_firstStep_partialProducts_compare_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:11]
  wire [8:0] quotient_secondGuess_firstStep_partialProducts_3 = {_quotient_secondGuess_firstStep_partialProducts_T_3
    , 3'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:22]
  wire [6:0] _GEN_22 = {{1'd0}, quotient_secondGuess_firstStep_partialProducts_0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 114:34]
  wire [7:0] _quotient_secondGuess_firstStep_partialSums_T = _GEN_22 + quotient_secondGuess_firstStep_partialProducts_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 114:34]
  wire [8:0] quotient_secondGuess_firstStep_partialSums_0 = _quotient_secondGuess_firstStep_partialSums_T +
    quotient_secondGuess_firstStep_partialProducts_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 114:39]
  wire [9:0] quotient_secondGuess_firstStep = quotient_secondGuess_firstStep_partialSums_0 +
    quotient_secondGuess_firstStep_partialProducts_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 111:15]
  wire  _quotient_secondGuess_firstStepRnd_roundedValue_T_4 = quotient_secondGuess_firstStep[2] & |
    quotient_secondGuess_firstStep[1:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 79:59]
  wire [5:0] _GEN_23 = {{5'd0}, _quotient_secondGuess_firstStepRnd_roundedValue_T_4}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 79:35]
  wire [6:0] quotient_secondGuess_firstStepRnd = quotient_secondGuess_firstStep[8:3] + _GEN_23; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 79:35]
  wire [5:0] _quotient_secondGuess_secondStep_T_1 = ~quotient_secondGuess_firstStepRnd[5:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 216:25]
  wire [5:0] quotient_secondGuess_secondStep = _quotient_secondGuess_secondStep_T_1 + 6'h1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 216:70]
  wire [5:0] quotient_secondGuess_finalStep_partialProducts_compare = quotient_secondGuess_secondStep[0] ? 6'h3f : 6'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 103:24]
  wire [5:0] quotient_secondGuess_finalStep_partialProducts_0 = quotient_initGuess &
    quotient_secondGuess_finalStep_partialProducts_compare; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:11]
  wire [5:0] quotient_secondGuess_finalStep_partialProducts_compare_1 = quotient_secondGuess_secondStep[1] ? 6'h3f : 6'h0
    ; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 103:24]
  wire [5:0] _quotient_secondGuess_finalStep_partialProducts_T_1 = quotient_initGuess &
    quotient_secondGuess_finalStep_partialProducts_compare_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:11]
  wire [6:0] quotient_secondGuess_finalStep_partialProducts_1 = {_quotient_secondGuess_finalStep_partialProducts_T_1
    , 1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:22]
  wire [5:0] quotient_secondGuess_finalStep_partialProducts_compare_2 = quotient_secondGuess_secondStep[2] ? 6'h3f : 6'h0
    ; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 103:24]
  wire [5:0] _quotient_secondGuess_finalStep_partialProducts_T_2 = quotient_initGuess &
    quotient_secondGuess_finalStep_partialProducts_compare_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:11]
  wire [7:0] quotient_secondGuess_finalStep_partialProducts_2 = {_quotient_secondGuess_finalStep_partialProducts_T_2
    , 2'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:22]
  wire [5:0] quotient_secondGuess_finalStep_partialProducts_compare_3 = quotient_secondGuess_secondStep[3] ? 6'h3f : 6'h0
    ; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 103:24]
  wire [5:0] _quotient_secondGuess_finalStep_partialProducts_T_3 = quotient_initGuess &
    quotient_secondGuess_finalStep_partialProducts_compare_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:11]
  wire [8:0] quotient_secondGuess_finalStep_partialProducts_3 = {_quotient_secondGuess_finalStep_partialProducts_T_3
    , 3'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:22]
  wire [5:0] quotient_secondGuess_finalStep_partialProducts_compare_4 = quotient_secondGuess_secondStep[4] ? 6'h3f : 6'h0
    ; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 103:24]
  wire [5:0] _quotient_secondGuess_finalStep_partialProducts_T_4 = quotient_initGuess &
    quotient_secondGuess_finalStep_partialProducts_compare_4; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:11]
  wire [9:0] quotient_secondGuess_finalStep_partialProducts_4 = {_quotient_secondGuess_finalStep_partialProducts_T_4
    , 4'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:22]
  wire [5:0] quotient_secondGuess_finalStep_partialProducts_compare_5 = quotient_secondGuess_secondStep[5] ? 6'h3f : 6'h0
    ; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 103:24]
  wire [5:0] _quotient_secondGuess_finalStep_partialProducts_T_5 = quotient_initGuess &
    quotient_secondGuess_finalStep_partialProducts_compare_5; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:11]
  wire [10:0] quotient_secondGuess_finalStep_partialProducts_5 = {_quotient_secondGuess_finalStep_partialProducts_T_5
    , 5'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:22]
  wire [6:0] _GEN_24 = {{1'd0}, quotient_secondGuess_finalStep_partialProducts_0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 114:34]
  wire [7:0] _quotient_secondGuess_finalStep_partialSums_T = _GEN_24 + quotient_secondGuess_finalStep_partialProducts_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 114:34]
  wire [8:0] quotient_secondGuess_finalStep_partialSums_0 = _quotient_secondGuess_finalStep_partialSums_T +
    quotient_secondGuess_finalStep_partialProducts_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 114:39]
  wire [9:0] _GEN_25 = {{1'd0}, quotient_secondGuess_finalStep_partialProducts_3}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 114:34]
  wire [10:0] _quotient_secondGuess_finalStep_partialSums_T_1 = _GEN_25 +
    quotient_secondGuess_finalStep_partialProducts_4; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 114:34]
  wire [11:0] quotient_secondGuess_finalStep_partialSums_1 = _quotient_secondGuess_finalStep_partialSums_T_1 +
    quotient_secondGuess_finalStep_partialProducts_5; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 114:39]
  wire [11:0] _GEN_26 = {{3'd0}, quotient_secondGuess_finalStep_partialSums_0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 111:15]
  wire [12:0] _quotient_secondGuess_finalStep_T = _GEN_26 + quotient_secondGuess_finalStep_partialSums_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 111:15]
  wire [11:0] quotient_secondGuess_finalStep = _quotient_secondGuess_finalStep_T[11:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 220:27 221:17]
  wire  _quotient_secondGuess_res_roundedValue_T_4 = quotient_secondGuess_finalStep[4] & |quotient_secondGuess_finalStep
    [3:2]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 79:59]
  wire [5:0] _GEN_27 = {{5'd0}, _quotient_secondGuess_res_roundedValue_T_4}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 79:35]
  wire [6:0] quotient_secondGuess = quotient_secondGuess_finalStep[10:5] + _GEN_27; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 79:35]
  wire [5:0] quotient_finalGuess_firstStep_partialProducts_0 = quotient_secondGuess[5:0] &
    quotient_secondGuess_firstStep_partialProducts_compare; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:11]
  wire [5:0] _quotient_finalGuess_firstStep_partialProducts_T_1 = quotient_secondGuess[5:0] &
    quotient_secondGuess_firstStep_partialProducts_compare_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:11]
  wire [6:0] quotient_finalGuess_firstStep_partialProducts_1 = {_quotient_finalGuess_firstStep_partialProducts_T_1
    , 1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:22]
  wire [5:0] _quotient_finalGuess_firstStep_partialProducts_T_2 = quotient_secondGuess[5:0] &
    quotient_secondGuess_firstStep_partialProducts_compare_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:11]
  wire [7:0] quotient_finalGuess_firstStep_partialProducts_2 = {_quotient_finalGuess_firstStep_partialProducts_T_2
    , 2'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:22]
  wire [5:0] _quotient_finalGuess_firstStep_partialProducts_T_3 = quotient_secondGuess[5:0] &
    quotient_secondGuess_firstStep_partialProducts_compare_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:11]
  wire [8:0] quotient_finalGuess_firstStep_partialProducts_3 = {_quotient_finalGuess_firstStep_partialProducts_T_3
    , 3'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:22]
  wire [6:0] _GEN_28 = {{1'd0}, quotient_finalGuess_firstStep_partialProducts_0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 114:34]
  wire [7:0] _quotient_finalGuess_firstStep_partialSums_T = _GEN_28 + quotient_finalGuess_firstStep_partialProducts_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 114:34]
  wire [8:0] quotient_finalGuess_firstStep_partialSums_0 = _quotient_finalGuess_firstStep_partialSums_T +
    quotient_finalGuess_firstStep_partialProducts_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 114:39]
  wire [9:0] quotient_finalGuess_firstStep = quotient_finalGuess_firstStep_partialSums_0 +
    quotient_finalGuess_firstStep_partialProducts_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 111:15]
  wire  _quotient_finalGuess_firstStepRnd_roundedValue_T_4 = quotient_finalGuess_firstStep[2] & |
    quotient_finalGuess_firstStep[1:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 79:59]
  wire [5:0] _GEN_29 = {{5'd0}, _quotient_finalGuess_firstStepRnd_roundedValue_T_4}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 79:35]
  wire [6:0] quotient_finalGuess_firstStepRnd = quotient_finalGuess_firstStep[8:3] + _GEN_29; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 79:35]
  wire [5:0] _quotient_finalGuess_secondStep_T_1 = ~quotient_finalGuess_firstStepRnd[5:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 216:25]
  wire [5:0] quotient_finalGuess_secondStep = _quotient_finalGuess_secondStep_T_1 + 6'h1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 216:70]
  wire [5:0] quotient_finalGuess_finalStep_partialProducts_compare = quotient_finalGuess_secondStep[0] ? 6'h3f : 6'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 103:24]
  wire [5:0] quotient_finalGuess_finalStep_partialProducts_0 = quotient_secondGuess[5:0] &
    quotient_finalGuess_finalStep_partialProducts_compare; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:11]
  wire [5:0] quotient_finalGuess_finalStep_partialProducts_compare_1 = quotient_finalGuess_secondStep[1] ? 6'h3f : 6'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 103:24]
  wire [5:0] _quotient_finalGuess_finalStep_partialProducts_T_1 = quotient_secondGuess[5:0] &
    quotient_finalGuess_finalStep_partialProducts_compare_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:11]
  wire [6:0] quotient_finalGuess_finalStep_partialProducts_1 = {_quotient_finalGuess_finalStep_partialProducts_T_1
    , 1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:22]
  wire [5:0] quotient_finalGuess_finalStep_partialProducts_compare_2 = quotient_finalGuess_secondStep[2] ? 6'h3f : 6'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 103:24]
  wire [5:0] _quotient_finalGuess_finalStep_partialProducts_T_2 = quotient_secondGuess[5:0] &
    quotient_finalGuess_finalStep_partialProducts_compare_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:11]
  wire [7:0] quotient_finalGuess_finalStep_partialProducts_2 = {_quotient_finalGuess_finalStep_partialProducts_T_2
    , 2'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:22]
  wire [5:0] quotient_finalGuess_finalStep_partialProducts_compare_3 = quotient_finalGuess_secondStep[3] ? 6'h3f : 6'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 103:24]
  wire [5:0] _quotient_finalGuess_finalStep_partialProducts_T_3 = quotient_secondGuess[5:0] &
    quotient_finalGuess_finalStep_partialProducts_compare_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:11]
  wire [8:0] quotient_finalGuess_finalStep_partialProducts_3 = {_quotient_finalGuess_finalStep_partialProducts_T_3
    , 3'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:22]
  wire [5:0] quotient_finalGuess_finalStep_partialProducts_compare_4 = quotient_finalGuess_secondStep[4] ? 6'h3f : 6'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 103:24]
  wire [5:0] _quotient_finalGuess_finalStep_partialProducts_T_4 = quotient_secondGuess[5:0] &
    quotient_finalGuess_finalStep_partialProducts_compare_4; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:11]
  wire [9:0] quotient_finalGuess_finalStep_partialProducts_4 = {_quotient_finalGuess_finalStep_partialProducts_T_4
    , 4'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:22]
  wire [5:0] quotient_finalGuess_finalStep_partialProducts_compare_5 = quotient_finalGuess_secondStep[5] ? 6'h3f : 6'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 103:24]
  wire [5:0] _quotient_finalGuess_finalStep_partialProducts_T_5 = quotient_secondGuess[5:0] &
    quotient_finalGuess_finalStep_partialProducts_compare_5; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:11]
  wire [10:0] quotient_finalGuess_finalStep_partialProducts_5 = {_quotient_finalGuess_finalStep_partialProducts_T_5
    , 5'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:22]
  wire [6:0] _GEN_30 = {{1'd0}, quotient_finalGuess_finalStep_partialProducts_0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 114:34]
  wire [7:0] _quotient_finalGuess_finalStep_partialSums_T = _GEN_30 + quotient_finalGuess_finalStep_partialProducts_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 114:34]
  wire [8:0] quotient_finalGuess_finalStep_partialSums_0 = _quotient_finalGuess_finalStep_partialSums_T +
    quotient_finalGuess_finalStep_partialProducts_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 114:39]
  wire [9:0] _GEN_31 = {{1'd0}, quotient_finalGuess_finalStep_partialProducts_3}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 114:34]
  wire [10:0] _quotient_finalGuess_finalStep_partialSums_T_1 = _GEN_31 + quotient_finalGuess_finalStep_partialProducts_4
    ; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 114:34]
  wire [11:0] quotient_finalGuess_finalStep_partialSums_1 = _quotient_finalGuess_finalStep_partialSums_T_1 +
    quotient_finalGuess_finalStep_partialProducts_5; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 114:39]
  wire [11:0] _GEN_32 = {{3'd0}, quotient_finalGuess_finalStep_partialSums_0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 111:15]
  wire [12:0] _quotient_finalGuess_finalStep_T = _GEN_32 + quotient_finalGuess_finalStep_partialSums_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 111:15]
  wire [11:0] quotient_finalGuess_finalStep = _quotient_finalGuess_finalStep_T[11:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 220:27 221:17]
  wire  _quotient_finalGuess_res_roundedValue_T_4 = quotient_finalGuess_finalStep[4] & |quotient_finalGuess_finalStep[3:
    2]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 79:59]
  wire [5:0] _GEN_33 = {{5'd0}, _quotient_finalGuess_res_roundedValue_T_4}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 79:35]
  wire [6:0] quotient_finalGuess = quotient_finalGuess_finalStep[10:5] + _GEN_33; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 79:35]
  wire [5:0] quotient_partialProducts_compare = dividendFraction[0] ? 6'h3f : 6'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 103:24]
  wire [5:0] quotient_partialProducts_0 = quotient_finalGuess[5:0] & quotient_partialProducts_compare; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:11]
  wire [5:0] quotient_partialProducts_compare_1 = dividendFraction[1] ? 6'h3f : 6'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 103:24]
  wire [5:0] _quotient_partialProducts_T_1 = quotient_finalGuess[5:0] & quotient_partialProducts_compare_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:11]
  wire [6:0] quotient_partialProducts_1 = {_quotient_partialProducts_T_1, 1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:22]
  wire [5:0] quotient_partialProducts_compare_2 = dividendFraction[2] ? 6'h3f : 6'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 103:24]
  wire [5:0] _quotient_partialProducts_T_2 = quotient_finalGuess[5:0] & quotient_partialProducts_compare_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:11]
  wire [7:0] quotient_partialProducts_2 = {_quotient_partialProducts_T_2, 2'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:22]
  wire [5:0] quotient_partialProducts_compare_3 = dividendFraction[3] ? 6'h3f : 6'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 103:24]
  wire [5:0] _quotient_partialProducts_T_3 = quotient_finalGuess[5:0] & quotient_partialProducts_compare_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:11]
  wire [8:0] quotient_partialProducts_3 = {_quotient_partialProducts_T_3, 3'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:22]
  wire [6:0] _GEN_34 = {{1'd0}, quotient_partialProducts_0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 114:34]
  wire [7:0] _quotient_partialSums_T = _GEN_34 + quotient_partialProducts_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 114:34]
  wire [8:0] quotient_partialSums_0 = _quotient_partialSums_T + quotient_partialProducts_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 114:39]
  wire [9:0] quotient = quotient_partialSums_0 + quotient_partialProducts_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 111:15]
  wire [7:0] _GEN_35 = {{4'd0}, quotient[7:4]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 60:44]
  wire [7:0] _leadingZeros_T_36 = _GEN_35 & 8'hf; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 60:44]
  wire [7:0] _leadingZeros_T_38 = {quotient[3:0], 4'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 60:44]
  wire [7:0] _leadingZeros_T_40 = _leadingZeros_T_38 & 8'hf0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 60:44]
  wire [7:0] _leadingZeros_T_41 = _leadingZeros_T_36 | _leadingZeros_T_40; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 60:44]
  wire [7:0] _GEN_36 = {{2'd0}, _leadingZeros_T_41[7:2]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 60:44]
  wire [7:0] _leadingZeros_T_46 = _GEN_36 & 8'h33; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 60:44]
  wire [7:0] _leadingZeros_T_48 = {_leadingZeros_T_41[5:0], 2'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 60:44]
  wire [7:0] _leadingZeros_T_50 = _leadingZeros_T_48 & 8'hcc; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 60:44]
  wire [7:0] _leadingZeros_T_51 = _leadingZeros_T_46 | _leadingZeros_T_50; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 60:44]
  wire [7:0] _GEN_37 = {{1'd0}, _leadingZeros_T_51[7:1]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 60:44]
  wire [7:0] _leadingZeros_T_56 = _GEN_37 & 8'h55; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 60:44]
  wire [7:0] _leadingZeros_T_58 = {_leadingZeros_T_51[6:0], 1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 60:44]
  wire [7:0] _leadingZeros_T_60 = _leadingZeros_T_58 & 8'haa; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 60:44]
  wire [7:0] _leadingZeros_T_61 = _leadingZeros_T_56 | _leadingZeros_T_60; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 60:44]
  wire [8:0] _leadingZeros_T_63 = {_leadingZeros_T_61,quotient[8]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 60:44]
  wire [3:0] _leadingZeros_T_73 = _leadingZeros_T_63[7] ? 4'h7 : 4'h8; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _leadingZeros_T_74 = _leadingZeros_T_63[6] ? 4'h6 : _leadingZeros_T_73; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _leadingZeros_T_75 = _leadingZeros_T_63[5] ? 4'h5 : _leadingZeros_T_74; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _leadingZeros_T_76 = _leadingZeros_T_63[4] ? 4'h4 : _leadingZeros_T_75; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _leadingZeros_T_77 = _leadingZeros_T_63[3] ? 4'h3 : _leadingZeros_T_76; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _leadingZeros_T_78 = _leadingZeros_T_63[2] ? 4'h2 : _leadingZeros_T_77; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _leadingZeros_T_79 = _leadingZeros_T_63[1] ? 4'h1 : _leadingZeros_T_78; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] shift = _leadingZeros_T_63[0] ? 4'h0 : _leadingZeros_T_79; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [9:0] _shiftedValue_T_33 = {quotient[8:0], 1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 65:23]
  wire [10:0] _shiftedValue_T_35 = {quotient[8:0], 2'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 65:23]
  wire [11:0] _shiftedValue_T_37 = {quotient[8:0], 3'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 65:23]
  wire [12:0] _shiftedValue_T_39 = {quotient[8:0], 4'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 65:23]
  wire [13:0] _shiftedValue_T_41 = {quotient[8:0], 5'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 65:23]
  wire [14:0] _shiftedValue_T_43 = {quotient[8:0], 6'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 65:23]
  wire [15:0] _shiftedValue_T_45 = {quotient[8:0], 7'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 65:23]
  wire [16:0] _shiftedValue_T_47 = {quotient[8:0], 8'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 65:23]
  wire [8:0] _shiftedValue_T_52 = 4'h1 == shift ? _shiftedValue_T_33[8:0] : quotient[8:0]; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [8:0] _shiftedValue_T_54 = 4'h2 == shift ? _shiftedValue_T_35[8:0] : _shiftedValue_T_52; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [8:0] _shiftedValue_T_56 = 4'h3 == shift ? _shiftedValue_T_37[8:0] : _shiftedValue_T_54; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [8:0] _shiftedValue_T_58 = 4'h4 == shift ? _shiftedValue_T_39[8:0] : _shiftedValue_T_56; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [8:0] _shiftedValue_T_60 = 4'h5 == shift ? _shiftedValue_T_41[8:0] : _shiftedValue_T_58; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [8:0] _shiftedValue_T_62 = 4'h6 == shift ? _shiftedValue_T_43[8:0] : _shiftedValue_T_60; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [8:0] _shiftedValue_T_64 = 4'h7 == shift ? _shiftedValue_T_45[8:0] : _shiftedValue_T_62; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [8:0] shiftedCalcValue = 4'h8 == shift ? _shiftedValue_T_47[8:0] : _shiftedValue_T_64; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [5:0] exponentShiftRight = 6'h0 - exponent_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 354:55]
  wire [5:0] exponentShiftLeft = exponent_1 - 6'h1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 357:35]
  wire  _T_2 = ~exponent_1[5]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 365:10]
  wire  _T_5 = ~exponent_1[5] & exponent_1[4:0] >= 5'hf; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 365:40]
  wire  _T_12 = _T_2 & exponent_1[4:0] < 5'hf; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 369:46]
  wire [4:0] _tempExponent_T_9 = exponent_1[4:0] + 5'h1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 371:51]
  wire  _tempFraction_T_2 = &quotient[1:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 375:59]
  wire [6:0] _GEN_38 = {{6'd0}, _tempFraction_T_2}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 374:81]
  wire [6:0] _tempFraction_T_4 = quotient[8:2] + _GEN_38; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 374:81]
  wire [4:0] _GEN_39 = {{1'd0}, shift}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 379:78]
  wire  _T_19 = _T_2 & exponent_1[4:0] > _GEN_39; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 379:46]
  wire [4:0] _tempExponent_T_12 = exponent_1[4:0] - _GEN_39; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 381:51]
  wire  _tempFraction_T_7 = &shiftedCalcValue[1:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 385:60]
  wire [6:0] _GEN_41 = {{6'd0}, _tempFraction_T_7}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 384:82]
  wire [6:0] _tempFraction_T_9 = shiftedCalcValue[8:2] + _GEN_41; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 384:82]
  wire [69:0] _GEN_0 = {{63'd0}, _tempFraction_T_4}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 395:74]
  wire [69:0] _tempFraction_T_15 = _GEN_0 << exponentShiftLeft; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 395:74]
  wire  _tempFraction_T_18 = &quotient[2:1]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 401:125]
  wire [6:0] _GEN_43 = {{6'd0}, _tempFraction_T_18}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 400:118]
  wire [6:0] _tempFraction_T_20 = quotient[9:3] + _GEN_43; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 400:118]
  wire [6:0] _tempFraction_T_21 = _tempFraction_T_20 >> exponentShiftRight; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 401:138]
  wire [69:0] _GEN_8 = _T_2 & exponent_1[4:0] > 5'h0 ? _tempFraction_T_15 : {{63'd0}, _tempFraction_T_21}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 391:82 392:22 400:22]
  wire [4:0] _GEN_9 = _T_19 & shiftedCalcValue[8] ? _tempExponent_T_12 : 5'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 380:55 381:20 390:20]
  wire [69:0] _GEN_10 = _T_19 & shiftedCalcValue[8] ? {{63'd0}, _tempFraction_T_9} : _GEN_8; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 380:55 382:20]
  wire [4:0] _GEN_11 = _T_12 & quotient[9] ? _tempExponent_T_9 : _GEN_9; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 370:54 371:20]
  wire [69:0] _GEN_12 = _T_12 & quotient[9] ? {{63'd0}, _tempFraction_T_4} : _GEN_10; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 370:54 372:20]
  wire [4:0] tempExponent_1 = _T_5 & quotient[9] ? 5'hf : _GEN_11; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 366:54 367:20]
  wire [69:0] _GEN_14 = _T_5 & quotient[9] ? 70'hff : _GEN_12; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 366:54 368:20]
  wire [7:0] tempFraction = _GEN_14[7:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 361:28]
  wire  _addOne_T_2 = roundingMode == 2'h0 & tempFraction[2]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 236:42]
  wire  _addOne_T_17 = _addOne_T_2 & ~tempFraction[1] & ~tempFraction[0] & tempFraction[3]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 237:90]
  wire  _addOne_T_18 = roundingMode == 2'h0 & tempFraction[2] & (tempFraction[1] | tempFraction[0]) | _addOne_T_17; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 236:102]
  wire  _addOne_T_24 = tempFraction[2] | tempFraction[1] | tempFraction[0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 238:70]
  wire  _addOne_T_27 = roundingMode == 2'h1 & (tempFraction[2] | tempFraction[1] | tempFraction[0]) & resultSign; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 238:90]
  wire  _addOne_T_28 = _addOne_T_18 | _addOne_T_27; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 237:110]
  wire  _addOne_T_38 = roundingMode == 2'h2 & _addOne_T_24 & ~resultSign; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 239:90]
  wire  addOne = _addOne_T_28 | _addOne_T_38; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 238:106]
  wire [3:0] _GEN_44 = {{3'd0}, addOne}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 241:66]
  wire [4:0] roundedFraction = tempFraction[6:3] + _GEN_44; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 241:66]
  wire [3:0] resultFraction = roundedFraction[4] ? roundedFraction[4:1] : roundedFraction[3:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 243:28]
  wire [4:0] _finalExponent_T_7 = tempExponent_1 + 5'h1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 247:20]
  wire [4:0] resultExponent = roundedFraction[4] | roundedFraction[3] & tempExponent_1 == 5'h0 ? _finalExponent_T_7 :
    tempExponent_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 246:28]
  wire  _overflow_T_9 = tempExponent_1 >= 5'hf & tempFraction[6:3] == 4'hf; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 252:42]
  wire  overflow = resultExponent > 5'hf | resultExponent[3:0] == 4'hf & resultFraction == 4'hf | _overflow_T_9; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 251:134]
  wire [4:0] resultStatus = {overflow,resultExponent == 5'h0,isResultNaN,1'h0,isResult0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 498:23]
  assign sign = enable & resultSign; // @[\\src\\main\\scala\\fpu8\\Divide.scala 23:24 24:10 30:10]
  assign exponent = enable ? resultExponent : 5'h0; // @[\\src\\main\\scala\\fpu8\\Divide.scala 23:24 25:14 31:14]
  assign fraction = enable ? resultFraction : 4'h0; // @[\\src\\main\\scala\\fpu8\\Divide.scala 23:24 26:14 32:14]
  assign status = enable ? resultStatus : 5'h0; // @[\\src\\main\\scala\\fpu8\\Divide.scala 23:24 27:12 33:12]
endmodule
module Compare(
  input        enable, // @[\\src\\main\\scala\\fpu8\\Compare.scala 6:18]
  input  [2:0] compareMode, // @[\\src\\main\\scala\\fpu8\\Compare.scala 7:23]
  input  [7:0] a_data, // @[\\src\\main\\scala\\fpu8\\Compare.scala 8:13]
  input  [7:0] b_data, // @[\\src\\main\\scala\\fpu8\\Compare.scala 9:13]
  output [7:0] z, // @[\\src\\main\\scala\\fpu8\\Compare.scala 10:13]
  output [4:0] status // @[\\src\\main\\scala\\fpu8\\Compare.scala 11:18]
);
  wire  _result_T_4 = a_data[6:3] == 4'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 35:39]
  wire  _result_T_6 = a_data[2:0] == 3'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 39:44]
  wire  _result_T_7 = _result_T_4 & _result_T_6; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 53:26]
  wire  _result_T_9 = b_data[6:3] == 4'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 35:39]
  wire  _result_T_11 = b_data[2:0] == 3'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 39:44]
  wire  _result_T_12 = _result_T_9 & _result_T_11; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 53:26]
  wire  _result_T_13 = _result_T_7 & _result_T_12; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 508:50]
  wire  _result_T_14 = ~(_result_T_7 & _result_T_12); // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 508:39]
  wire  _result_T_20 = a_data[6:0] > b_data[6:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 29:77]
  wire  _result_T_21 = a_data[7] & _result_T_20; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 509:26]
  wire  _result_T_22 = a_data[7] > b_data[7] & ~(_result_T_7 & _result_T_12) | _result_T_21; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 508:65]
  wire  _result_T_24 = ~a_data[7]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 509:67]
  wire  _result_T_27 = a_data[6:0] < b_data[6:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 31:74]
  wire [7:0] result_result = _result_T_22 | ~a_data[7] & _result_T_27 ? 8'h38 : 8'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 509:99 511:14 513:14]
  wire  _result_T_51 = a_data[7] & _result_T_27; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 523:26]
  wire  _result_T_52 = a_data[7] < b_data[7] & _result_T_14 | _result_T_51; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 522:65]
  wire [7:0] result_result_1 = _result_T_52 | _result_T_24 & _result_T_20 ? 8'h38 : 8'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 523:100 525:14 527:14]
  wire [7:0] result_result_2 = a_data == b_data | _result_T_13 ? 8'h38 : 8'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 536:65 538:14 540:14]
  wire [7:0] _result_T_116 = result_result ^ result_result_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 548:20]
  wire [7:0] _result_T_160 = result_result_1 ^ result_result_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 554:20]
  wire  _T_6 = compareMode == 3'h5; // @[\\src\\main\\scala\\fpu8\\Compare.scala 28:28]
  wire  _result_T_176 = a_data[6:3] == 4'hf; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 37:41]
  wire  _result_T_178 = a_data[2:0] == 3'h7; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 41:46]
  wire  _result_T_179 = _result_T_176 & _result_T_178; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 43:30]
  wire  _result_T_181 = b_data[6:3] == 4'hf; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 37:41]
  wire  _result_T_183 = b_data[2:0] == 3'h7; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 41:46]
  wire  _result_T_184 = _result_T_181 & _result_T_183; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 43:30]
  wire [7:0] result_result_7 = a_data != b_data & _result_T_14 | _result_T_179 & _result_T_184 ? 8'h38 : 8'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 561:99 563:14 565:14]
  wire [7:0] _GEN_8 = compareMode == 3'h5 ? result_result_7 : 8'h0; // @[\\src\\main\\scala\\fpu8\\Compare.scala 28:36 29:14 31:14]
  wire [7:0] _GEN_9 = compareMode == 3'h4 ? _result_T_160 : _GEN_8; // @[\\src\\main\\scala\\fpu8\\Compare.scala 26:37 27:14]
  wire [7:0] _GEN_10 = compareMode == 3'h3 ? _result_T_116 : _GEN_9; // @[\\src\\main\\scala\\fpu8\\Compare.scala 24:37 25:14]
  wire [7:0] _GEN_11 = compareMode == 3'h2 ? result_result_2 : _GEN_10; // @[\\src\\main\\scala\\fpu8\\Compare.scala 22:37 23:14]
  wire [7:0] _GEN_12 = compareMode == 3'h1 ? result_result_1 : _GEN_11; // @[\\src\\main\\scala\\fpu8\\Compare.scala 20:37 21:14]
  wire [7:0] _GEN_13 = compareMode == 3'h0 ? result_result : _GEN_12; // @[\\src\\main\\scala\\fpu8\\Compare.scala 18:31 19:14]
  wire [7:0] result = enable ? _GEN_13 : 8'h0; // @[\\src\\main\\scala\\fpu8\\Compare.scala 17:23 48:12]
  wire [7:0] _z_T_13 = _T_6 & _result_T_179 & _result_T_184 ? result : 8'h0; // @[\\src\\main\\scala\\fpu8\\Compare.scala 39:15]
  wire  is0 = enable & _result_T_13; // @[\\src\\main\\scala\\fpu8\\Compare.scala 17:23 35:9 51:9]
  wire  isNaN = enable & (_result_T_179 | _result_T_184); // @[\\src\\main\\scala\\fpu8\\Compare.scala 17:23 34:11 50:11]
  wire [2:0] _GEN_16 = isNaN ? 3'h4 : {{2'd0}, is0}; // @[\\src\\main\\scala\\fpu8\\Compare.scala 37:16 38:14]
  wire [7:0] _GEN_17 = isNaN ? _z_T_13 : result; // @[\\src\\main\\scala\\fpu8\\Compare.scala 37:16 39:9]
  wire [2:0] _GEN_21 = enable ? _GEN_16 : 3'h0; // @[\\src\\main\\scala\\fpu8\\Compare.scala 17:23 52:12]
  assign z = enable ? _GEN_17 : 8'h0; // @[\\src\\main\\scala\\fpu8\\Compare.scala 17:23 49:7]
  assign status = {{2'd0}, _GEN_21};
endmodule
module Convert(
  input        enable, // @[\\src\\main\\scala\\fpu8\\Convert.scala 6:18]
  input  [7:0] a_data, // @[\\src\\main\\scala\\fpu8\\Convert.scala 7:13]
  output [7:0] z, // @[\\src\\main\\scala\\fpu8\\Convert.scala 10:13]
  output [4:0] status // @[\\src\\main\\scala\\fpu8\\Convert.scala 11:18]
);
  wire  _fraction_T_1 = a_data[6:3] == 4'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 35:39]
  wire  _fraction_T_2 = ~_fraction_T_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 572:24]
  wire [3:0] fraction = {_fraction_T_2,a_data[2:0]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 572:23]
  wire [3:0] _leadingZeros_T_8 = {fraction[0],fraction[1],fraction[2],fraction[3]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 60:44]
  wire [1:0] _leadingZeros_T_13 = _leadingZeros_T_8[2] ? 2'h2 : 2'h3; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [1:0] _leadingZeros_T_14 = _leadingZeros_T_8[1] ? 2'h1 : _leadingZeros_T_13; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [1:0] shift = _leadingZeros_T_8[0] ? 2'h0 : _leadingZeros_T_14; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [4:0] _shiftedValue_T_3 = {fraction, 1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 65:23]
  wire [5:0] _shiftedValue_T_5 = {fraction, 2'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 65:23]
  wire [6:0] _shiftedValue_T_7 = {fraction, 3'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 65:23]
  wire [3:0] _shiftedValue_T_10 = 2'h1 == shift ? _shiftedValue_T_3[3:0] : fraction; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [3:0] _shiftedValue_T_12 = 2'h2 == shift ? _shiftedValue_T_5[3:0] : _shiftedValue_T_10; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [3:0] shiftedFraction = 2'h3 == shift ? _shiftedValue_T_7[3:0] : _shiftedValue_T_12; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [3:0] _GEN_8 = {{2'd0}, shift}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 575:40]
  wire [4:0] _tempExponent_T_2 = 4'h9 - _GEN_8; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 575:40]
  wire [4:0] _tempExponent_T_5 = 4'h8 + a_data[6:3]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 575:54]
  wire [4:0] tempExponent = _fraction_T_1 ? _tempExponent_T_2 : _tempExponent_T_5; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 575:27]
  wire [2:0] tempFraction = shiftedFraction[3:1]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 576:39]
  wire  addOne = |a_data[6:3] & &shiftedFraction[1:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 578:38]
  wire [2:0] _GEN_9 = {{2'd0}, addOne}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 580:40]
  wire [3:0] roundedFraction = tempFraction + _GEN_9; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 580:40]
  wire [4:0] _finalExponent_T_3 = tempExponent + 5'h1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 582:83]
  wire [4:0] finalExponent = roundedFraction[3] ? _finalExponent_T_3 : tempExponent; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 582:28]
  wire [2:0] finalFraction = roundedFraction[3] ? roundedFraction[3:1] : roundedFraction[2:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 583:28]
  wire  _T_4 = a_data[2:0] == 3'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 39:44]
  wire  _T_5 = _fraction_T_1 & _T_4; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 53:26]
  wire  _T_8 = a_data[6:3] == 4'hf; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 37:41]
  wire  _T_10 = a_data[2:0] == 3'h7; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 41:46]
  wire  _T_11 = _T_8 & _T_10; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 43:30]
  wire  _T_12 = ~_T_11; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 590:18]
  wire [7:0] _result_T_2 = {a_data[7],finalExponent,finalFraction[1:0]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 591:20]
  wire [7:0] _result_T_4 = {a_data[7],5'h0,2'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 594:20]
  wire [7:0] _GEN_0 = _T_11 ? 8'h7f : 8'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 596:23 597:14 600:14]
  wire [2:0] _GEN_1 = _T_11 ? 3'h4 : 3'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 596:23 598:14 601:14]
  wire [7:0] _GEN_2 = _T_5 & _T_12 ? _result_T_4 : _GEN_0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 593:31 594:14]
  wire [2:0] _GEN_3 = _T_5 & _T_12 ? 3'h1 : _GEN_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 593:31 595:14]
  wire [7:0] result = ~_T_5 & ~_T_11 ? _result_T_2 : _GEN_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 590:26 591:14]
  wire [2:0] _GEN_5 = ~_T_5 & ~_T_11 ? 3'h0 : _GEN_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 590:26 592:14]
  wire [4:0] resultStatus = {{2'd0}, _GEN_5}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 588:22]
  assign z = enable ? result : 8'h0; // @[\\src\\main\\scala\\fpu8\\Convert.scala 13:23 19:7 22:7]
  assign status = enable ? resultStatus : 5'h0; // @[\\src\\main\\scala\\fpu8\\Convert.scala 13:23 20:12 23:12]
endmodule
module GenerateFinalResult(
  input        enable, // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 12:18]
  input        sign, // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 13:16]
  input  [3:0] exponent, // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 14:20]
  input  [2:0] mantissa, // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 15:20]
  input  [1:0] roundingMode, // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 16:24]
  input        overflow, // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 17:20]
  input        saturationMode, // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 18:26]
  input        is0, // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 20:15]
  input        isNaN, // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 21:17]
  output [7:0] z // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 23:13]
);
  wire  _result_T_4 = ~isNaN; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 40:18]
  wire  _result_T_6 = roundingMode == 2'h0; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 42:28]
  wire  _result_T_7 = ~saturationMode; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 42:54]
  wire  _result_T_9 = roundingMode == 2'h1; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 43:26]
  wire  _result_T_10 = roundingMode == 2'h2; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 43:50]
  wire  _result_T_14 = ~sign; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 43:93]
  wire  _result_T_15 = (roundingMode == 2'h1 | roundingMode == 2'h2) & _result_T_7 & ~sign; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 43:85]
  wire  _result_T_16 = roundingMode == 2'h0 & ~saturationMode | _result_T_15; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 42:63]
  wire [7:0] _result_z_T_1 = {sign,4'hf,3'h6}; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 46:19]
  wire [7:0] _GEN_0 = _result_T_9 & sign | _result_T_10 & saturationMode & _result_T_14 ? 8'h7e : 8'h0; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 49:128 50:13 52:13]
  wire [7:0] _GEN_1 = _result_T_9 & saturationMode & _result_T_14 | _result_T_10 & sign ? 8'hfe : _GEN_0; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 47:128 48:13]
  wire [7:0] _GEN_2 = _result_T_6 & saturationMode | roundingMode == 2'h3 & _result_T_7 ? _result_z_T_1 : _GEN_1; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 45:122 46:13]
  wire [7:0] _GEN_3 = _result_T_16 ? 8'h7f : _GEN_2; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 43:103 44:13]
  wire [7:0] _result_z_T_4 = {sign,exponent,mantissa}; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 55:17]
  wire [7:0] _GEN_4 = overflow ? _GEN_3 : _result_z_T_4; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 41:22 55:11]
  wire [7:0] _GEN_5 = isNaN ? 8'h7f : 8'h0; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 59:23 60:9 62:9]
  wire [7:0] _GEN_6 = is0 & _result_T_4 ? 8'h0 : _GEN_5; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 57:31 58:9]
  wire [7:0] result = ~is0 & ~isNaN ? _GEN_4 : _GEN_6; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 40:26]
  assign z = enable ? result : 8'h0; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 31:23 32:7 34:7]
endmodule
module FPU8Generator(
  input        clock,
  input        reset,
  input        enable, // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 9:18]
  input  [7:0] a_data, // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 10:13]
  input  [7:0] b_data, // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 11:13]
  input  [3:0] opCode, // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 12:18]
  input  [1:0] roundingMode, // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 13:24]
  input        saturationMode, // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 14:26]
  output [7:0] z, // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 15:13]
  output [4:0] status // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 16:18]
);
  wire  addSub_enable; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 18:22]
  wire [7:0] addSub_a_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 18:22]
  wire [7:0] addSub_b_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 18:22]
  wire  addSub_subtract; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 18:22]
  wire [1:0] addSub_roundingMode; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 18:22]
  wire  addSub_sign; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 18:22]
  wire [4:0] addSub_exponent; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 18:22]
  wire [3:0] addSub_fraction; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 18:22]
  wire [4:0] addSub_status; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 18:22]
  wire  multiply_enable; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 20:24]
  wire [7:0] multiply_a_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 20:24]
  wire [7:0] multiply_b_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 20:24]
  wire [1:0] multiply_roundingMode; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 20:24]
  wire  multiply_sign; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 20:24]
  wire [4:0] multiply_exponent; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 20:24]
  wire [3:0] multiply_fraction; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 20:24]
  wire [4:0] multiply_status; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 20:24]
  wire  divide_enable; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 22:22]
  wire [7:0] divide_a_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 22:22]
  wire [7:0] divide_b_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 22:22]
  wire [1:0] divide_roundingMode; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 22:22]
  wire  divide_sign; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 22:22]
  wire [4:0] divide_exponent; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 22:22]
  wire [3:0] divide_fraction; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 22:22]
  wire [4:0] divide_status; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 22:22]
  wire  compare_enable; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 24:23]
  wire [2:0] compare_compareMode; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 24:23]
  wire [7:0] compare_a_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 24:23]
  wire [7:0] compare_b_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 24:23]
  wire [7:0] compare_z; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 24:23]
  wire [4:0] compare_status; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 24:23]
  wire  convert_enable; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 26:23]
  wire [7:0] convert_a_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 26:23]
  wire [7:0] convert_z; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 26:23]
  wire [4:0] convert_status; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 26:23]
  wire  generateFinalResult_enable; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 28:35]
  wire  generateFinalResult_sign; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 28:35]
  wire [3:0] generateFinalResult_exponent; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 28:35]
  wire [2:0] generateFinalResult_mantissa; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 28:35]
  wire [1:0] generateFinalResult_roundingMode; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 28:35]
  wire  generateFinalResult_overflow; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 28:35]
  wire  generateFinalResult_saturationMode; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 28:35]
  wire  generateFinalResult_is0; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 28:35]
  wire  generateFinalResult_isNaN; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 28:35]
  wire [7:0] generateFinalResult_z; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 28:35]
  wire  _addSub_enable_T_2 = opCode == 4'h0 | opCode == 4'h1; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 30:39]
  wire  _multiply_enable_T = opCode == 4'h2; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 36:33]
  wire  _divide_enable_T = opCode == 4'h3; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 41:31]
  wire  _compare_enable_T = opCode == 4'h4; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 46:32]
  wire  _compare_enable_T_1 = opCode == 4'h5; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 46:50]
  wire  _compare_enable_T_3 = opCode == 4'h6; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 46:68]
  wire  _compare_enable_T_5 = opCode == 4'h7; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 46:86]
  wire  _compare_enable_T_7 = opCode == 4'h8; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 46:104]
  wire  _compare_enable_T_10 = opCode == 4'h4 | opCode == 4'h5 | opCode == 4'h6 | opCode == 4'h7 | opCode == 4'h8 |
    opCode == 4'h9; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 46:112]
  wire [2:0] _compare_compareMode_T_5 = _compare_enable_T_7 ? 3'h4 : 3'h5; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 52:14]
  wire [2:0] _compare_compareMode_T_6 = _compare_enable_T_5 ? 3'h3 : _compare_compareMode_T_5; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 51:12]
  wire [2:0] _compare_compareMode_T_7 = _compare_enable_T_3 ? 3'h2 : _compare_compareMode_T_6; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 50:10]
  wire [2:0] _compare_compareMode_T_8 = _compare_enable_T_1 ? 3'h1 : _compare_compareMode_T_7; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 49:8]
  wire  _convert_enable_T = opCode == 4'ha; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 56:32]
  wire [7:0] _GEN_1 = _convert_enable_T ? convert_z : 8'h0; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 119:30 131:7 145:7]
  wire [4:0] _GEN_2 = _convert_enable_T ? convert_status : 5'h0; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 119:30 132:12 146:12]
  wire [7:0] _GEN_4 = _compare_enable_T_10 ? compare_z : _GEN_1; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 105:119 117:7]
  wire [4:0] _GEN_5 = _compare_enable_T_10 ? compare_status : _GEN_2; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 105:119 118:12]
  wire  _GEN_6 = _divide_enable_T & divide_sign; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 91:30 92:30]
  wire [3:0] _GEN_7 = _divide_enable_T ? divide_exponent[3:0] : 4'h0; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 91:30 93:34]
  wire [2:0] _GEN_8 = _divide_enable_T ? divide_fraction[2:0] : 3'h0; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 91:30 94:34]
  wire [1:0] _GEN_9 = _divide_enable_T ? roundingMode : 2'h0; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 91:30 95:38]
  wire  _GEN_10 = _divide_enable_T & divide_status[4]; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 91:30 96:34]
  wire  _GEN_11 = _divide_enable_T & saturationMode; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 91:30 97:40]
  wire  _GEN_13 = _divide_enable_T & divide_status[0]; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 91:30 99:29]
  wire  _GEN_14 = _divide_enable_T & divide_status[2]; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 91:30 100:31]
  wire [7:0] _GEN_16 = _divide_enable_T ? generateFinalResult_z : _GEN_4; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 91:30 103:7]
  wire [4:0] _GEN_17 = _divide_enable_T ? divide_status : _GEN_5; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 104:12 91:30]
  wire  _GEN_18 = _multiply_enable_T ? multiply_sign : _GEN_6; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 77:30 78:30]
  wire [3:0] _GEN_19 = _multiply_enable_T ? multiply_exponent[3:0] : _GEN_7; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 77:30 79:34]
  wire [2:0] _GEN_20 = _multiply_enable_T ? multiply_fraction[2:0] : _GEN_8; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 77:30 80:34]
  wire [1:0] _GEN_21 = _multiply_enable_T ? roundingMode : _GEN_9; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 77:30 81:38]
  wire  _GEN_22 = _multiply_enable_T ? multiply_status[4] : _GEN_10; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 77:30 82:34]
  wire  _GEN_23 = _multiply_enable_T ? saturationMode : _GEN_11; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 77:30 83:40]
  wire  _GEN_25 = _multiply_enable_T ? multiply_status[0] : _GEN_13; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 77:30 85:29]
  wire  _GEN_26 = _multiply_enable_T ? multiply_status[2] : _GEN_14; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 77:30 86:31]
  wire [7:0] _GEN_28 = _multiply_enable_T ? generateFinalResult_z : _GEN_16; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 77:30 89:7]
  wire [4:0] _GEN_29 = _multiply_enable_T ? multiply_status : _GEN_17; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 77:30 90:12]
  Add addSub ( // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 18:22]
    .enable(addSub_enable),
    .a_data(addSub_a_data),
    .b_data(addSub_b_data),
    .subtract(addSub_subtract),
    .roundingMode(addSub_roundingMode),
    .sign(addSub_sign),
    .exponent(addSub_exponent),
    .fraction(addSub_fraction),
    .status(addSub_status)
  );
  Multiply multiply ( // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 20:24]
    .enable(multiply_enable),
    .a_data(multiply_a_data),
    .b_data(multiply_b_data),
    .roundingMode(multiply_roundingMode),
    .sign(multiply_sign),
    .exponent(multiply_exponent),
    .fraction(multiply_fraction),
    .status(multiply_status)
  );
  Divide divide ( // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 22:22]
    .enable(divide_enable),
    .a_data(divide_a_data),
    .b_data(divide_b_data),
    .roundingMode(divide_roundingMode),
    .sign(divide_sign),
    .exponent(divide_exponent),
    .fraction(divide_fraction),
    .status(divide_status)
  );
  Compare compare ( // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 24:23]
    .enable(compare_enable),
    .compareMode(compare_compareMode),
    .a_data(compare_a_data),
    .b_data(compare_b_data),
    .z(compare_z),
    .status(compare_status)
  );
  Convert convert ( // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 26:23]
    .enable(convert_enable),
    .a_data(convert_a_data),
    .z(convert_z),
    .status(convert_status)
  );
  GenerateFinalResult generateFinalResult ( // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 28:35]
    .enable(generateFinalResult_enable),
    .sign(generateFinalResult_sign),
    .exponent(generateFinalResult_exponent),
    .mantissa(generateFinalResult_mantissa),
    .roundingMode(generateFinalResult_roundingMode),
    .overflow(generateFinalResult_overflow),
    .saturationMode(generateFinalResult_saturationMode),
    .is0(generateFinalResult_is0),
    .isNaN(generateFinalResult_isNaN),
    .z(generateFinalResult_z)
  );
  assign z = _addSub_enable_T_2 ? generateFinalResult_z : _GEN_28; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 63:42 75:7]
  assign status = _addSub_enable_T_2 ? addSub_status : _GEN_29; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 63:42 76:12]
  assign addSub_enable = (opCode == 4'h0 | opCode == 4'h1) & enable; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 30:23]
  assign addSub_a_data = a_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 31:12]
  assign addSub_b_data = b_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 32:12]
  assign addSub_subtract = opCode == 4'h1; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 33:33]
  assign addSub_roundingMode = roundingMode; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 34:23]
  assign multiply_enable = opCode == 4'h2 & enable; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 36:25]
  assign multiply_a_data = a_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 37:14]
  assign multiply_b_data = b_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 38:14]
  assign multiply_roundingMode = roundingMode; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 39:25]
  assign divide_enable = opCode == 4'h3 & enable; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 41:23]
  assign divide_a_data = a_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 42:12]
  assign divide_b_data = b_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 43:12]
  assign divide_roundingMode = roundingMode; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 44:23]
  assign compare_enable = (opCode == 4'h4 | opCode == 4'h5 | opCode == 4'h6 | opCode == 4'h7 | opCode == 4'h8 | opCode
     == 4'h9) & enable; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 46:24]
  assign compare_compareMode = _compare_enable_T ? 3'h0 : _compare_compareMode_T_8; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 48:29]
  assign compare_a_data = a_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 53:13]
  assign compare_b_data = b_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 54:13]
  assign convert_enable = opCode == 4'ha & enable; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 56:24]
  assign convert_a_data = a_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 57:13]
  assign generateFinalResult_enable = enable; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 61:30]
  assign generateFinalResult_sign = _addSub_enable_T_2 ? addSub_sign : _GEN_18; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 63:42 64:30]
  assign generateFinalResult_exponent = _addSub_enable_T_2 ? addSub_exponent[3:0] : _GEN_19; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 63:42 65:34]
  assign generateFinalResult_mantissa = _addSub_enable_T_2 ? addSub_fraction[2:0] : _GEN_20; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 63:42 66:34]
  assign generateFinalResult_roundingMode = _addSub_enable_T_2 ? roundingMode : _GEN_21; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 63:42 67:38]
  assign generateFinalResult_overflow = _addSub_enable_T_2 ? addSub_status[4] : _GEN_22; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 63:42 68:34]
  assign generateFinalResult_saturationMode = _addSub_enable_T_2 ? saturationMode : _GEN_23; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 63:42 69:40]
  assign generateFinalResult_is0 = _addSub_enable_T_2 ? addSub_status[0] : _GEN_25; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 63:42 71:29]
  assign generateFinalResult_isNaN = _addSub_enable_T_2 ? addSub_status[2] : _GEN_26; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 63:42 72:31]
endmodule
