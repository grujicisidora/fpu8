module Add(
  input        enable, // @[\\src\\main\\scala\\fpu8\\Add.scala 9:18]
  input  [7:0] a_data, // @[\\src\\main\\scala\\fpu8\\Add.scala 10:13]
  input  [7:0] b_data, // @[\\src\\main\\scala\\fpu8\\Add.scala 11:13]
  input        subtract, // @[\\src\\main\\scala\\fpu8\\Add.scala 12:20]
  input  [1:0] roundingMode, // @[\\src\\main\\scala\\fpu8\\Add.scala 13:24]
  output       sign, // @[\\src\\main\\scala\\fpu8\\Add.scala 14:16]
  output [5:0] exponent, // @[\\src\\main\\scala\\fpu8\\Add.scala 15:20]
  output [2:0] fraction, // @[\\src\\main\\scala\\fpu8\\Add.scala 16:20]
  output       overflow, // @[\\src\\main\\scala\\fpu8\\Add.scala 17:20]
  output       isInfty, // @[\\src\\main\\scala\\fpu8\\Add.scala 18:19]
  output       is0, // @[\\src\\main\\scala\\fpu8\\Add.scala 19:15]
  output       isNaN, // @[\\src\\main\\scala\\fpu8\\Add.scala 20:17]
  output       NaNFractionValue // @[\\src\\main\\scala\\fpu8\\Add.scala 21:28]
);
  wire  compare = a_data[6:0] > b_data[6:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 29:77]
  wire [7:0] greaterOperand_data = compare ? a_data : b_data; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 124:29]
  wire [7:0] smallerOperand_data = compare ? b_data : a_data; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 125:29]
  wire  resultSign = compare ? a_data[7] : b_data[7] ^ subtract; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 126:19]
  wire  subtraction = subtract ^ greaterOperand_data[7] ^ smallerOperand_data[7]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 127:54]
  wire [4:0] exponent_1 = greaterOperand_data[6:2]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 25:28]
  wire  _greaterOperandFraction_T_1 = exponent_1 == 5'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 33:39]
  wire  _greaterOperandFraction_T_2 = ~_greaterOperandFraction_T_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 129:38]
  wire  _smallerOperandFraction_T_1 = smallerOperand_data[6:2] == 5'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 33:39]
  wire  _smallerOperandFraction_T_2 = ~_smallerOperandFraction_T_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 130:38]
  wire  isOnlySmallerDenormalized = _greaterOperandFraction_T_2 & _smallerOperandFraction_T_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 131:60]
  wire [4:0] _shift_T_2 = exponent_1 - 5'h1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 134:31]
  wire [4:0] _shift_T_6 = exponent_1 - smallerOperand_data[6:2]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 135:31]
  wire [4:0] shift = isOnlySmallerDenormalized ? _shift_T_2 : _shift_T_6; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 132:20]
  wire  _shiftedFraction_shifted_T = shift >= 5'h5; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 140:15]
  wire [7:0] _shiftedFraction_shifted_T_1 = {5'h0,_smallerOperandFraction_T_2,smallerOperand_data[1:0]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 141:12]
  wire [7:0] _shiftedFraction_shifted_T_2 = {_smallerOperandFraction_T_2,smallerOperand_data[1:0],5'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 142:12]
  wire [7:0] _shiftedFraction_shifted_T_3 = _shiftedFraction_shifted_T_2 >> shift; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 142:54]
  wire [7:0] shiftedFraction_shifted = _shiftedFraction_shifted_T ? _shiftedFraction_shifted_T_1 :
    _shiftedFraction_shifted_T_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 139:24]
  wire [5:0] smallerOperandFraction_1 = {shiftedFraction_shifted[7:3],|shiftedFraction_shifted[2:0]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 144:10]
  wire [5:0] greaterOperandFraction_1 = {_greaterOperandFraction_T_2,greaterOperand_data[1:0],3'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 146:45]
  wire  _isResultNaN_T_1 = a_data[6:2] == 5'h1f; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 35:41]
  wire  _isResultNaN_T_3 = a_data[1:0] == 2'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 37:44]
  wire  _isResultNaN_T_4 = ~_isResultNaN_T_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 42:15]
  wire  _isResultNaN_T_5 = _isResultNaN_T_1 & _isResultNaN_T_4; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 41:30]
  wire  _isResultNaN_T_7 = b_data[6:2] == 5'h1f; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 35:41]
  wire  _isResultNaN_T_9 = b_data[1:0] == 2'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 37:44]
  wire  _isResultNaN_T_10 = ~_isResultNaN_T_9; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 42:15]
  wire  _isResultNaN_T_11 = _isResultNaN_T_7 & _isResultNaN_T_10; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 41:30]
  wire  _isResultNaN_T_17 = _isResultNaN_T_1 & _isResultNaN_T_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 47:24]
  wire  _isResultNaN_T_22 = _isResultNaN_T_7 & _isResultNaN_T_9; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 47:24]
  wire  isResultNaN = _isResultNaN_T_5 | _isResultNaN_T_11 | _isResultNaN_T_17 & _isResultNaN_T_22 & subtraction; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 392:57]
  wire  _isResultInfty_T_11 = ~isResultNaN; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 397:65]
  wire  isResultInfty = (_isResultNaN_T_17 | _isResultNaN_T_22) & ~isResultNaN; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 397:63]
  wire  _isResult0_T_2 = a_data[6:0] == b_data[6:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 31:77]
  wire  isResult0 = _isResult0_T_2 & subtraction & _isResultInfty_T_11 & ~isResultInfty; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 401:101]
  wire  resultNaNFractionValue = a_data[1:0] > b_data[1:0] ? a_data[0] : b_data[0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 118:18]
  wire [6:0] _calculatedValue_T_1 = greaterOperandFraction_1 - smallerOperandFraction_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 406:32]
  wire [6:0] _calculatedValue_T_3 = greaterOperandFraction_1 + smallerOperandFraction_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 407:32]
  wire [6:0] calculatedValue = subtraction ? _calculatedValue_T_1 : _calculatedValue_T_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 405:32]
  wire [7:0] paddedCalcValue = {calculatedValue,1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 262:15]
  wire [6:0] _leadingZeros_T_17 = {paddedCalcValue[0],paddedCalcValue[1],paddedCalcValue[2],paddedCalcValue[3],
    paddedCalcValue[4],paddedCalcValue[5],paddedCalcValue[6]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 58:44]
  wire [2:0] _leadingZeros_T_25 = _leadingZeros_T_17[5] ? 3'h5 : 3'h6; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] _leadingZeros_T_26 = _leadingZeros_T_17[4] ? 3'h4 : _leadingZeros_T_25; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] _leadingZeros_T_27 = _leadingZeros_T_17[3] ? 3'h3 : _leadingZeros_T_26; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] _leadingZeros_T_28 = _leadingZeros_T_17[2] ? 3'h2 : _leadingZeros_T_27; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] _leadingZeros_T_29 = _leadingZeros_T_17[1] ? 3'h1 : _leadingZeros_T_28; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] shift_1 = _leadingZeros_T_17[0] ? 3'h0 : _leadingZeros_T_29; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [13:0] _GEN_5 = {{7'd0}, paddedCalcValue[6:0]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 60:27]
  wire [13:0] _shiftedValue_T = _GEN_5 << shift_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 60:27]
  wire  _T_1 = &exponent_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 270:19]
  wire [4:0] _tempExponent_T_1 = exponent_1 + 5'h1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 274:32]
  wire [6:0] _tempFraction_T_3 = {paddedCalcValue[7:2],|paddedCalcValue[1:0]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 275:26]
  wire [4:0] _GEN_15 = {{2'd0}, shift_1}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 276:25]
  wire [6:0] shiftedCalcValue = _shiftedValue_T[6:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 56:28 60:18]
  wire [4:0] _tempExponent_T_3 = exponent_1 - _GEN_15; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 277:32]
  wire [37:0] _GEN_7 = {{31'd0}, paddedCalcValue[6:0]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 282:47]
  wire [37:0] _tempFraction_T_7 = _GEN_7 << _shift_T_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 282:47]
  wire [37:0] _GEN_0 = exponent_1 > 5'h0 ? _tempFraction_T_7 : {{31'd0}, paddedCalcValue[6:0]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 281:28 282:22 284:22]
  wire [4:0] _GEN_1 = exponent_1 > _GEN_15 & shiftedCalcValue[6] ? _tempExponent_T_3 : 5'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 276:57 277:20 280:20]
  wire [37:0] _GEN_2 = exponent_1 > _GEN_15 & shiftedCalcValue[6] ? {{31'd0}, shiftedCalcValue} : _GEN_0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 276:57 278:20]
  wire [4:0] _GEN_3 = ~_T_1 & paddedCalcValue[7] ? _tempExponent_T_1 : _GEN_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 273:54 274:20]
  wire [37:0] _GEN_4 = ~_T_1 & paddedCalcValue[7] ? {{31'd0}, _tempFraction_T_3} : _GEN_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 273:54 275:20]
  wire [4:0] tempExponent = &exponent_1 & paddedCalcValue[7] ? exponent_1 : _GEN_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 270:47 271:20]
  wire [37:0] _GEN_6 = &exponent_1 & paddedCalcValue[7] ? 38'h7f : _GEN_4; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 270:47 272:20]
  wire [6:0] tempFraction = _GEN_6[6:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 268:28]
  wire  _addOne_T_2 = roundingMode == 2'h0 & tempFraction[3]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 229:42]
  wire  _addOne_T_17 = _addOne_T_2 & ~tempFraction[2] & ~tempFraction[1] & tempFraction[4]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 230:90]
  wire  _addOne_T_18 = roundingMode == 2'h0 & tempFraction[3] & (tempFraction[2] | tempFraction[1]) | _addOne_T_17; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 229:102]
  wire  _addOne_T_24 = tempFraction[3] | tempFraction[2] | tempFraction[1]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 231:70]
  wire  _addOne_T_27 = roundingMode == 2'h1 & (tempFraction[3] | tempFraction[2] | tempFraction[1]) & resultSign; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 231:90]
  wire  _addOne_T_28 = _addOne_T_18 | _addOne_T_27; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 230:110]
  wire  _addOne_T_38 = roundingMode == 2'h2 & _addOne_T_24 & ~resultSign; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 232:90]
  wire  addOne = _addOne_T_28 | _addOne_T_38; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 231:106]
  wire [2:0] _GEN_17 = {{2'd0}, addOne}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 234:66]
  wire [3:0] roundedFraction = tempFraction[6:4] + _GEN_17; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 234:66]
  wire [2:0] resultFraction = roundedFraction[3] ? roundedFraction[3:1] : roundedFraction[2:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 236:28]
  wire [4:0] _finalExponent_T_7 = tempExponent + 5'h1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 240:20]
  wire [4:0] resultExponent = roundedFraction[3] | roundedFraction[2] & tempExponent == 5'h0 ? _finalExponent_T_7 :
    tempExponent; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 239:28]
  wire  resultOverflow = tempExponent == 5'h1f; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 243:76]
  wire [4:0] _GEN_8 = enable ? resultExponent : 5'h0; // @[\\src\\main\\scala\\fpu8\\Add.scala 26:24 28:14 37:14]
  assign sign = enable & resultSign; // @[\\src\\main\\scala\\fpu8\\Add.scala 26:24 27:10 36:10]
  assign exponent = {{1'd0}, _GEN_8};
  assign fraction = enable ? resultFraction : 3'h0; // @[\\src\\main\\scala\\fpu8\\Add.scala 26:24 29:14 38:14]
  assign overflow = enable & resultOverflow; // @[\\src\\main\\scala\\fpu8\\Add.scala 26:24 30:14 39:14]
  assign isInfty = enable & isResultInfty; // @[\\src\\main\\scala\\fpu8\\Add.scala 26:24 31:13 40:13]
  assign is0 = enable & isResult0; // @[\\src\\main\\scala\\fpu8\\Add.scala 26:24 32:9 41:9]
  assign isNaN = enable & isResultNaN; // @[\\src\\main\\scala\\fpu8\\Add.scala 26:24 33:11 42:11]
  assign NaNFractionValue = enable & resultNaNFractionValue; // @[\\src\\main\\scala\\fpu8\\Add.scala 26:24 34:22 43:22]
endmodule
module Multiply(
  input        enable, // @[\\src\\main\\scala\\fpu8\\Multiply.scala 9:18]
  input  [7:0] a_data, // @[\\src\\main\\scala\\fpu8\\Multiply.scala 10:13]
  input  [7:0] b_data, // @[\\src\\main\\scala\\fpu8\\Multiply.scala 11:13]
  input  [1:0] roundingMode, // @[\\src\\main\\scala\\fpu8\\Multiply.scala 12:24]
  output       sign, // @[\\src\\main\\scala\\fpu8\\Multiply.scala 13:16]
  output [5:0] exponent, // @[\\src\\main\\scala\\fpu8\\Multiply.scala 14:20]
  output [2:0] fraction, // @[\\src\\main\\scala\\fpu8\\Multiply.scala 15:20]
  output       overflow, // @[\\src\\main\\scala\\fpu8\\Multiply.scala 16:20]
  output       isInfty, // @[\\src\\main\\scala\\fpu8\\Multiply.scala 17:19]
  output       is0, // @[\\src\\main\\scala\\fpu8\\Multiply.scala 18:15]
  output       isNaN, // @[\\src\\main\\scala\\fpu8\\Multiply.scala 19:17]
  output       NaNFractionValue // @[\\src\\main\\scala\\fpu8\\Multiply.scala 20:28]
);
  wire  _isResultNaN_T_1 = a_data[6:2] == 5'h1f; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 35:41]
  wire  _isResultNaN_T_3 = a_data[1:0] == 2'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 37:44]
  wire  _isResultNaN_T_4 = _isResultNaN_T_1 & _isResultNaN_T_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 47:24]
  wire  _isResultNaN_T_6 = b_data[6:2] == 5'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 33:39]
  wire  _isResultNaN_T_8 = b_data[1:0] == 2'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 37:44]
  wire  _isResultNaN_T_9 = _isResultNaN_T_6 & _isResultNaN_T_8; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 51:26]
  wire  _isResultNaN_T_15 = ~_isResultNaN_T_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 42:15]
  wire  _isResultNaN_T_16 = _isResultNaN_T_1 & _isResultNaN_T_15; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 41:30]
  wire  _isResultNaN_T_19 = b_data[6:2] == 5'h1f; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 35:41]
  wire  _isResultNaN_T_22 = _isResultNaN_T_19 & _isResultNaN_T_8; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 47:24]
  wire  _isResultNaN_T_24 = a_data[6:2] == 5'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 33:39]
  wire  _isResultNaN_T_27 = _isResultNaN_T_24 & _isResultNaN_T_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 51:26]
  wire  _isResultNaN_T_34 = ~_isResultNaN_T_8; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 42:15]
  wire  _isResultNaN_T_35 = _isResultNaN_T_19 & _isResultNaN_T_34; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 41:30]
  wire  isResultNaN = _isResultNaN_T_4 & _isResultNaN_T_9 | _isResultNaN_T_16 | _isResultNaN_T_22 & _isResultNaN_T_27 |
    _isResultNaN_T_35; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 420:104]
  wire  _isResultInfty_T_18 = ~_isResultNaN_T_35; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 425:62]
  wire  _isResultInfty_T_38 = ~_isResultNaN_T_16; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 425:110]
  wire  isResultInfty = _isResultNaN_T_4 & ~_isResultNaN_T_9 & ~_isResultNaN_T_35 | _isResultNaN_T_22 & ~
    _isResultNaN_T_27 & ~_isResultNaN_T_16; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 425:76]
  wire  isResult0 = _isResultNaN_T_27 & _isResultInfty_T_18 | _isResultNaN_T_9 & _isResultInfty_T_38; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 429:62]
  wire  resultNaNFractionValue = a_data[1:0] > b_data[1:0] ? a_data[0] : b_data[0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 118:18]
  wire  resultSign = a_data[7] ^ b_data[7]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 151:26]
  wire [6:0] _exponent_T_11 = {2'h0,a_data[6:2]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 163:16]
  wire [6:0] _exponent_T_13 = {2'h0,b_data[6:2]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 163:47]
  wire [6:0] _exponent_T_15 = _exponent_T_11 + _exponent_T_13; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 163:42]
  wire [6:0] _exponent_T_17 = _exponent_T_15 - 7'he; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 163:74]
  wire [6:0] _exponent_T_25 = _exponent_T_15 - 7'hf; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 164:74]
  wire [6:0] _exponent_T_26 = _isResultNaN_T_24 ^ _isResultNaN_T_6 ? _exponent_T_17 : _exponent_T_25; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 162:14]
  wire [6:0] exponent_1 = _isResultNaN_T_24 & _isResultNaN_T_6 ? 7'h1c : _exponent_T_26; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 160:12]
  wire  _firstOperandFraction_T_2 = ~_isResultNaN_T_24; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 166:36]
  wire [2:0] firstOperandFraction = {_firstOperandFraction_T_2,a_data[1:0]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 166:35]
  wire  _secondOperandFraction_T_2 = ~_isResultNaN_T_6; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 167:37]
  wire [2:0] secondOperandFraction = {_secondOperandFraction_T_2,b_data[1:0]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 167:36]
  wire [2:0] product_partialProducts_compare = secondOperandFraction[0] ? 3'h7 : 3'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 96:24]
  wire [2:0] product_partialProducts_0 = firstOperandFraction & product_partialProducts_compare; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 97:11]
  wire [2:0] product_partialProducts_compare_1 = secondOperandFraction[1] ? 3'h7 : 3'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 96:24]
  wire [2:0] _product_partialProducts_T_1 = firstOperandFraction & product_partialProducts_compare_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 97:11]
  wire [3:0] product_partialProducts_1 = {_product_partialProducts_T_1, 1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 97:22]
  wire [2:0] product_partialProducts_compare_2 = secondOperandFraction[2] ? 3'h7 : 3'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 96:24]
  wire [2:0] _product_partialProducts_T_2 = firstOperandFraction & product_partialProducts_compare_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 97:11]
  wire [4:0] product_partialProducts_2 = {_product_partialProducts_T_2, 2'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 97:22]
  wire [3:0] _GEN_15 = {{1'd0}, product_partialProducts_0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 107:34]
  wire [4:0] _product_partialSums_T = _GEN_15 + product_partialProducts_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 107:34]
  wire [5:0] product = _product_partialSums_T + product_partialProducts_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 107:39]
  wire [4:0] _leadingZeros_T_11 = {product[0],product[1],product[2],product[3],product[4]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 58:44]
  wire [2:0] _leadingZeros_T_17 = _leadingZeros_T_11[3] ? 3'h3 : 3'h4; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] _leadingZeros_T_18 = _leadingZeros_T_11[2] ? 3'h2 : _leadingZeros_T_17; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] _leadingZeros_T_19 = _leadingZeros_T_11[1] ? 3'h1 : _leadingZeros_T_18; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] shift = _leadingZeros_T_11[0] ? 3'h0 : _leadingZeros_T_19; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [11:0] _GEN_7 = {{7'd0}, product[4:0]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 60:27]
  wire [11:0] _shiftedValue_T = _GEN_7 << shift; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 60:27]
  wire [6:0] exponentShiftRight = 7'h0 - exponent_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 296:58]
  wire [6:0] exponentShiftLeft = exponent_1 - 7'h1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 298:38]
  wire  _T_2 = ~exponent_1[6]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 304:10]
  wire  _T_5 = ~exponent_1[6] & exponent_1[5:0] >= 6'h1f; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 304:40]
  wire  _T_12 = _T_2 & exponent_1[5:0] < 6'h1f; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 308:46]
  wire [4:0] _tempExponent_T_2 = exponent_1[4:0] + 5'h1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 310:38]
  wire [4:0] _tempFraction_T_3 = {product[5:2],|product[1:0]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 311:26]
  wire [5:0] _GEN_16 = {{3'd0}, shift}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 312:78]
  wire  _T_19 = _T_2 & exponent_1[5:0] > _GEN_16; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 312:46]
  wire [4:0] shiftedCalcValue = _shiftedValue_T[4:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 56:28 60:18]
  wire [5:0] _tempExponent_T_5 = exponent_1[5:0] - _GEN_16; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 314:51]
  wire [131:0] _GEN_9 = {{127'd0}, product[4:0]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 319:71]
  wire [131:0] _tempFraction_T_5 = _GEN_9 << exponentShiftLeft; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 319:71]
  wire [4:0] _tempFraction_T_10 = _tempFraction_T_3 >> exponentShiftRight; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 321:110]
  wire [131:0] _GEN_0 = _T_2 & exponent_1[5:0] > 6'h0 ? _tempFraction_T_5 : {{127'd0}, _tempFraction_T_10}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 318:82 319:22 321:22]
  wire [5:0] _GEN_1 = _T_19 & shiftedCalcValue[4] ? _tempExponent_T_5 : 6'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 313:55 314:20 317:20]
  wire [131:0] _GEN_2 = _T_19 & shiftedCalcValue[4] ? {{127'd0}, shiftedCalcValue} : _GEN_0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 313:55 315:20]
  wire [5:0] _GEN_3 = _T_12 & product[5] ? {{1'd0}, _tempExponent_T_2} : _GEN_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 309:54 310:20]
  wire [131:0] _GEN_4 = _T_12 & product[5] ? {{127'd0}, _tempFraction_T_3} : _GEN_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 309:54 311:20]
  wire [5:0] _GEN_5 = _T_5 & product[5] ? 6'h1f : _GEN_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 305:54 306:20]
  wire [131:0] _GEN_6 = _T_5 & product[5] ? 132'h1f : _GEN_4; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 305:54 307:20]
  wire [4:0] tempFraction = _GEN_6[4:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 302:28]
  wire  _addOne_T_2 = roundingMode == 2'h0 & tempFraction[2]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 229:42]
  wire  _addOne_T_17 = _addOne_T_2 & ~tempFraction[1] & ~tempFraction[0] & tempFraction[3]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 230:90]
  wire  _addOne_T_18 = roundingMode == 2'h0 & tempFraction[2] & (tempFraction[1] | tempFraction[0]) | _addOne_T_17; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 229:102]
  wire  _addOne_T_24 = tempFraction[2] | tempFraction[1] | tempFraction[0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 231:70]
  wire  _addOne_T_27 = roundingMode == 2'h1 & (tempFraction[2] | tempFraction[1] | tempFraction[0]) & resultSign; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 231:90]
  wire  _addOne_T_28 = _addOne_T_18 | _addOne_T_27; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 230:110]
  wire  _addOne_T_38 = roundingMode == 2'h2 & _addOne_T_24 & ~resultSign; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 232:90]
  wire  addOne = _addOne_T_28 | _addOne_T_38; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 231:106]
  wire [2:0] _GEN_18 = {{2'd0}, addOne}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 234:66]
  wire [3:0] roundedFraction = tempFraction[4:2] + _GEN_18; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 234:66]
  wire [2:0] resultFraction = roundedFraction[3] ? roundedFraction[3:1] : roundedFraction[2:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 236:28]
  wire [4:0] tempExponent = _GEN_5[4:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 300:28]
  wire [4:0] _finalExponent_T_7 = tempExponent + 5'h1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 240:20]
  wire [4:0] resultExponent = roundedFraction[3] | roundedFraction[2] & tempExponent == 5'h0 ? _finalExponent_T_7 :
    tempExponent; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 239:28]
  wire  resultOverflow = tempExponent == 5'h1f; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 243:76]
  wire [4:0] _GEN_8 = enable ? resultExponent : 5'h0; // @[\\src\\main\\scala\\fpu8\\Multiply.scala 25:24 27:14 36:14]
  assign sign = enable & resultSign; // @[\\src\\main\\scala\\fpu8\\Multiply.scala 25:24 26:10 35:10]
  assign exponent = {{1'd0}, _GEN_8};
  assign fraction = enable ? resultFraction : 3'h0; // @[\\src\\main\\scala\\fpu8\\Multiply.scala 25:24 28:14 37:14]
  assign overflow = enable & resultOverflow; // @[\\src\\main\\scala\\fpu8\\Multiply.scala 25:24 29:14 38:14]
  assign isInfty = enable & isResultInfty; // @[\\src\\main\\scala\\fpu8\\Multiply.scala 25:24 30:13 39:13]
  assign is0 = enable & isResult0; // @[\\src\\main\\scala\\fpu8\\Multiply.scala 25:24 31:9 40:9]
  assign isNaN = enable & isResultNaN; // @[\\src\\main\\scala\\fpu8\\Multiply.scala 25:24 32:11 41:11]
  assign NaNFractionValue = enable & resultNaNFractionValue; // @[\\src\\main\\scala\\fpu8\\Multiply.scala 25:24 33:22 42:22]
endmodule
module Divide(
  input        enable, // @[\\src\\main\\scala\\fpu8\\Divide.scala 9:18]
  input  [7:0] a_data, // @[\\src\\main\\scala\\fpu8\\Divide.scala 10:13]
  input  [7:0] b_data, // @[\\src\\main\\scala\\fpu8\\Divide.scala 11:13]
  input  [1:0] roundingMode, // @[\\src\\main\\scala\\fpu8\\Divide.scala 12:24]
  output       sign, // @[\\src\\main\\scala\\fpu8\\Divide.scala 13:16]
  output [5:0] exponent, // @[\\src\\main\\scala\\fpu8\\Divide.scala 14:20]
  output [2:0] fraction, // @[\\src\\main\\scala\\fpu8\\Divide.scala 15:20]
  output       overflow, // @[\\src\\main\\scala\\fpu8\\Divide.scala 16:20]
  output       isInfty, // @[\\src\\main\\scala\\fpu8\\Divide.scala 17:19]
  output       is0, // @[\\src\\main\\scala\\fpu8\\Divide.scala 18:15]
  output       isNaN, // @[\\src\\main\\scala\\fpu8\\Divide.scala 19:17]
  output       NaNFractionValue // @[\\src\\main\\scala\\fpu8\\Divide.scala 20:28]
);
  wire  _isResultNaN_T_1 = a_data[6:2] == 5'h1f; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 35:41]
  wire  _isResultNaN_T_3 = a_data[1:0] == 2'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 37:44]
  wire  _isResultNaN_T_4 = ~_isResultNaN_T_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 42:15]
  wire  _isResultNaN_T_5 = _isResultNaN_T_1 & _isResultNaN_T_4; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 41:30]
  wire  _isResultNaN_T_7 = b_data[6:2] == 5'h1f; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 35:41]
  wire  _isResultNaN_T_9 = b_data[1:0] == 2'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 37:44]
  wire  _isResultNaN_T_10 = ~_isResultNaN_T_9; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 42:15]
  wire  _isResultNaN_T_11 = _isResultNaN_T_7 & _isResultNaN_T_10; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 41:30]
  wire  _isResultNaN_T_14 = a_data[6:2] == 5'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 33:39]
  wire  _isResultNaN_T_17 = _isResultNaN_T_14 & _isResultNaN_T_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 51:26]
  wire  _isResultNaN_T_19 = b_data[6:2] == 5'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 33:39]
  wire  _isResultNaN_T_22 = _isResultNaN_T_19 & _isResultNaN_T_9; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 51:26]
  wire  _isResultNaN_T_29 = _isResultNaN_T_1 & _isResultNaN_T_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 47:24]
  wire  _isResultNaN_T_34 = _isResultNaN_T_7 & _isResultNaN_T_9; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 47:24]
  wire  isResultNaN = _isResultNaN_T_5 | _isResultNaN_T_11 | _isResultNaN_T_17 & _isResultNaN_T_22 | _isResultNaN_T_29
     & _isResultNaN_T_34; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 448:84]
  wire  _isResultInfty_T_17 = ~_isResultNaN_T_29; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 453:58]
  wire  _isResultInfty_T_25 = ~_isResultNaN_T_5; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 453:75]
  wire  _isResultInfty_T_38 = ~_isResultNaN_T_11; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 453:108]
  wire  isResultInfty = _isResultNaN_T_22 & ~_isResultNaN_T_17 & ~_isResultNaN_T_29 & ~_isResultNaN_T_5 |
    _isResultNaN_T_29 & ~_isResultNaN_T_11; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 453:88]
  wire  isResult0 = _isResultNaN_T_17 & ~_isResultNaN_T_22 & _isResultInfty_T_38 | _isResultNaN_T_34 &
    _isResultInfty_T_17 & _isResultInfty_T_25; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 458:72]
  wire  resultNaNFractionValue = a_data[1:0] > b_data[1:0] ? a_data[0] : b_data[0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 118:18]
  wire  resultSign = a_data[7] ^ b_data[7]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 173:26]
  wire [2:0] _tempDividendFraction_T_3 = {a_data[1:0],1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 175:10]
  wire [2:0] _tempDividendFraction_T_5 = {1'h1,a_data[1:0]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 176:10]
  wire [2:0] tempDividendFraction = _isResultNaN_T_14 ? _tempDividendFraction_T_3 : _tempDividendFraction_T_5; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 174:35]
  wire [2:0] _tempDivisorFraction_T_3 = {b_data[1:0],1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 179:10]
  wire [2:0] _tempDivisorFraction_T_5 = {1'h1,b_data[1:0]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 180:10]
  wire [2:0] tempDivisorFraction = _isResultNaN_T_19 ? _tempDivisorFraction_T_3 : _tempDivisorFraction_T_5; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 178:34]
  wire [6:0] _tempExponent_T_1 = {2'h0,a_data[6:2]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 182:27]
  wire [6:0] _tempExponent_T_3 = {2'h0,b_data[6:2]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 183:10]
  wire [6:0] _tempExponent_T_5 = _tempExponent_T_1 - _tempExponent_T_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 182:53]
  wire [6:0] tempExponent = _tempExponent_T_5 + 7'hf; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 183:37]
  wire [2:0] _leadingZeros_T_5 = {tempDividendFraction[0],tempDividendFraction[1],tempDividendFraction[2]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 58:44]
  wire [1:0] _leadingZeros_T_9 = _leadingZeros_T_5[1] ? 2'h1 : 2'h2; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [1:0] dividendShift = _leadingZeros_T_5[0] ? 2'h0 : _leadingZeros_T_9; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _GEN_0 = {{3'd0}, tempDividendFraction}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 60:27]
  wire [5:0] _shiftedValue_T = _GEN_0 << dividendShift; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 60:27]
  wire [2:0] _leadingZeros_T_16 = {tempDivisorFraction[0],tempDivisorFraction[1],tempDivisorFraction[2]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 58:44]
  wire [1:0] _leadingZeros_T_20 = _leadingZeros_T_16[1] ? 2'h1 : 2'h2; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [1:0] divisorShift = _leadingZeros_T_16[0] ? 2'h0 : _leadingZeros_T_20; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _GEN_9 = {{3'd0}, tempDivisorFraction}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 60:27]
  wire [5:0] _shiftedValue_T_1 = _GEN_9 << divisorShift; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 60:27]
  wire [6:0] _GEN_19 = {{5'd0}, dividendShift}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 190:33]
  wire [6:0] _exponent_T_1 = tempExponent - _GEN_19; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 190:33]
  wire [6:0] _GEN_20 = {{5'd0}, divisorShift}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 190:49]
  wire [6:0] exponent_1 = _exponent_T_1 + _GEN_20; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 190:49]
  wire [2:0] divisorFraction = _shiftedValue_T_1[2:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 56:28 60:18]
  wire [2:0] _GEN_1 = 2'h1 == divisorFraction[1:0] ? 3'h5 : 3'h7; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 198:{24,24}]
  wire [2:0] _GEN_2 = 2'h2 == divisorFraction[1:0] ? 3'h3 : _GEN_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 198:{24,24}]
  wire [2:0] _GEN_3 = 2'h3 == divisorFraction[1:0] ? 3'h1 : _GEN_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 198:{24,24}]
  wire [4:0] quotient_initGuess = {2'h1,_GEN_3}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 198:24]
  wire [4:0] quotient_secondGuess_firstStep_partialProducts_compare = divisorFraction[0] ? 5'h1f : 5'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 96:24]
  wire [4:0] quotient_secondGuess_firstStep_partialProducts_0 = quotient_initGuess &
    quotient_secondGuess_firstStep_partialProducts_compare; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 97:11]
  wire [4:0] quotient_secondGuess_firstStep_partialProducts_compare_1 = divisorFraction[1] ? 5'h1f : 5'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 96:24]
  wire [4:0] _quotient_secondGuess_firstStep_partialProducts_T_1 = quotient_initGuess &
    quotient_secondGuess_firstStep_partialProducts_compare_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 97:11]
  wire [5:0] quotient_secondGuess_firstStep_partialProducts_1 = {_quotient_secondGuess_firstStep_partialProducts_T_1
    , 1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 97:22]
  wire [4:0] quotient_secondGuess_firstStep_partialProducts_compare_2 = divisorFraction[2] ? 5'h1f : 5'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 96:24]
  wire [4:0] _quotient_secondGuess_firstStep_partialProducts_T_2 = quotient_initGuess &
    quotient_secondGuess_firstStep_partialProducts_compare_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 97:11]
  wire [6:0] quotient_secondGuess_firstStep_partialProducts_2 = {_quotient_secondGuess_firstStep_partialProducts_T_2
    , 2'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 97:22]
  wire [5:0] _GEN_21 = {{1'd0}, quotient_secondGuess_firstStep_partialProducts_0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 107:34]
  wire [6:0] _quotient_secondGuess_firstStep_partialSums_T = _GEN_21 + quotient_secondGuess_firstStep_partialProducts_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 107:34]
  wire [7:0] quotient_secondGuess_firstStep = _quotient_secondGuess_firstStep_partialSums_T +
    quotient_secondGuess_firstStep_partialProducts_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 107:39]
  wire [5:0] quotient_secondGuess_firstStepRnd = {1'h0,quotient_secondGuess_firstStep[6:2]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 74:12]
  wire [4:0] _quotient_secondGuess_secondStep_T_1 = ~quotient_secondGuess_firstStepRnd[4:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 209:25]
  wire [4:0] quotient_secondGuess_secondStep = _quotient_secondGuess_secondStep_T_1 + 5'h1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 209:70]
  wire [4:0] quotient_secondGuess_finalStep_partialProducts_compare = quotient_secondGuess_secondStep[0] ? 5'h1f : 5'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 96:24]
  wire [4:0] quotient_secondGuess_finalStep_partialProducts_0 = quotient_initGuess &
    quotient_secondGuess_finalStep_partialProducts_compare; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 97:11]
  wire [4:0] quotient_secondGuess_finalStep_partialProducts_compare_1 = quotient_secondGuess_secondStep[1] ? 5'h1f : 5'h0
    ; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 96:24]
  wire [4:0] _quotient_secondGuess_finalStep_partialProducts_T_1 = quotient_initGuess &
    quotient_secondGuess_finalStep_partialProducts_compare_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 97:11]
  wire [5:0] quotient_secondGuess_finalStep_partialProducts_1 = {_quotient_secondGuess_finalStep_partialProducts_T_1
    , 1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 97:22]
  wire [4:0] quotient_secondGuess_finalStep_partialProducts_compare_2 = quotient_secondGuess_secondStep[2] ? 5'h1f : 5'h0
    ; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 96:24]
  wire [4:0] _quotient_secondGuess_finalStep_partialProducts_T_2 = quotient_initGuess &
    quotient_secondGuess_finalStep_partialProducts_compare_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 97:11]
  wire [6:0] quotient_secondGuess_finalStep_partialProducts_2 = {_quotient_secondGuess_finalStep_partialProducts_T_2
    , 2'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 97:22]
  wire [4:0] quotient_secondGuess_finalStep_partialProducts_compare_3 = quotient_secondGuess_secondStep[3] ? 5'h1f : 5'h0
    ; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 96:24]
  wire [4:0] _quotient_secondGuess_finalStep_partialProducts_T_3 = quotient_initGuess &
    quotient_secondGuess_finalStep_partialProducts_compare_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 97:11]
  wire [7:0] quotient_secondGuess_finalStep_partialProducts_3 = {_quotient_secondGuess_finalStep_partialProducts_T_3
    , 3'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 97:22]
  wire [4:0] quotient_secondGuess_finalStep_partialProducts_compare_4 = quotient_secondGuess_secondStep[4] ? 5'h1f : 5'h0
    ; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 96:24]
  wire [4:0] _quotient_secondGuess_finalStep_partialProducts_T_4 = quotient_initGuess &
    quotient_secondGuess_finalStep_partialProducts_compare_4; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 97:11]
  wire [8:0] quotient_secondGuess_finalStep_partialProducts_4 = {_quotient_secondGuess_finalStep_partialProducts_T_4
    , 4'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 97:22]
  wire [5:0] _GEN_22 = {{1'd0}, quotient_secondGuess_finalStep_partialProducts_0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 107:34]
  wire [6:0] _quotient_secondGuess_finalStep_partialSums_T = _GEN_22 + quotient_secondGuess_finalStep_partialProducts_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 107:34]
  wire [7:0] quotient_secondGuess_finalStep_partialSums_0 = _quotient_secondGuess_finalStep_partialSums_T +
    quotient_secondGuess_finalStep_partialProducts_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 107:39]
  wire [8:0] _GEN_23 = {{1'd0}, quotient_secondGuess_finalStep_partialProducts_3}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 108:31]
  wire [9:0] quotient_secondGuess_finalStep_partialSums_1 = _GEN_23 + quotient_secondGuess_finalStep_partialProducts_4; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 108:31]
  wire [9:0] _GEN_24 = {{2'd0}, quotient_secondGuess_finalStep_partialSums_0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:15]
  wire [10:0] _quotient_secondGuess_finalStep_T = _GEN_24 + quotient_secondGuess_finalStep_partialSums_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:15]
  wire [9:0] quotient_secondGuess_finalStep = _quotient_secondGuess_finalStep_T[9:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 213:27 214:17]
  wire  _quotient_secondGuess_res_roundedValue_T_4 = quotient_secondGuess_finalStep[3] & |quotient_secondGuess_finalStep
    [2:1]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 72:59]
  wire [4:0] _GEN_25 = {{4'd0}, _quotient_secondGuess_res_roundedValue_T_4}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 72:35]
  wire [5:0] quotient_secondGuess = quotient_secondGuess_finalStep[8:4] + _GEN_25; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 72:35]
  wire [4:0] quotient_finalGuess_firstStep_partialProducts_0 = quotient_secondGuess[4:0] &
    quotient_secondGuess_firstStep_partialProducts_compare; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 97:11]
  wire [4:0] _quotient_finalGuess_firstStep_partialProducts_T_1 = quotient_secondGuess[4:0] &
    quotient_secondGuess_firstStep_partialProducts_compare_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 97:11]
  wire [5:0] quotient_finalGuess_firstStep_partialProducts_1 = {_quotient_finalGuess_firstStep_partialProducts_T_1
    , 1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 97:22]
  wire [4:0] _quotient_finalGuess_firstStep_partialProducts_T_2 = quotient_secondGuess[4:0] &
    quotient_secondGuess_firstStep_partialProducts_compare_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 97:11]
  wire [6:0] quotient_finalGuess_firstStep_partialProducts_2 = {_quotient_finalGuess_firstStep_partialProducts_T_2
    , 2'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 97:22]
  wire [5:0] _GEN_26 = {{1'd0}, quotient_finalGuess_firstStep_partialProducts_0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 107:34]
  wire [6:0] _quotient_finalGuess_firstStep_partialSums_T = _GEN_26 + quotient_finalGuess_firstStep_partialProducts_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 107:34]
  wire [7:0] quotient_finalGuess_firstStep = _quotient_finalGuess_firstStep_partialSums_T +
    quotient_finalGuess_firstStep_partialProducts_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 107:39]
  wire [5:0] quotient_finalGuess_firstStepRnd = {1'h0,quotient_finalGuess_firstStep[6:2]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 74:12]
  wire [4:0] _quotient_finalGuess_secondStep_T_1 = ~quotient_finalGuess_firstStepRnd[4:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 209:25]
  wire [4:0] quotient_finalGuess_secondStep = _quotient_finalGuess_secondStep_T_1 + 5'h1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 209:70]
  wire [4:0] quotient_finalGuess_finalStep_partialProducts_compare = quotient_finalGuess_secondStep[0] ? 5'h1f : 5'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 96:24]
  wire [4:0] quotient_finalGuess_finalStep_partialProducts_0 = quotient_secondGuess[4:0] &
    quotient_finalGuess_finalStep_partialProducts_compare; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 97:11]
  wire [4:0] quotient_finalGuess_finalStep_partialProducts_compare_1 = quotient_finalGuess_secondStep[1] ? 5'h1f : 5'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 96:24]
  wire [4:0] _quotient_finalGuess_finalStep_partialProducts_T_1 = quotient_secondGuess[4:0] &
    quotient_finalGuess_finalStep_partialProducts_compare_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 97:11]
  wire [5:0] quotient_finalGuess_finalStep_partialProducts_1 = {_quotient_finalGuess_finalStep_partialProducts_T_1
    , 1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 97:22]
  wire [4:0] quotient_finalGuess_finalStep_partialProducts_compare_2 = quotient_finalGuess_secondStep[2] ? 5'h1f : 5'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 96:24]
  wire [4:0] _quotient_finalGuess_finalStep_partialProducts_T_2 = quotient_secondGuess[4:0] &
    quotient_finalGuess_finalStep_partialProducts_compare_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 97:11]
  wire [6:0] quotient_finalGuess_finalStep_partialProducts_2 = {_quotient_finalGuess_finalStep_partialProducts_T_2
    , 2'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 97:22]
  wire [4:0] quotient_finalGuess_finalStep_partialProducts_compare_3 = quotient_finalGuess_secondStep[3] ? 5'h1f : 5'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 96:24]
  wire [4:0] _quotient_finalGuess_finalStep_partialProducts_T_3 = quotient_secondGuess[4:0] &
    quotient_finalGuess_finalStep_partialProducts_compare_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 97:11]
  wire [7:0] quotient_finalGuess_finalStep_partialProducts_3 = {_quotient_finalGuess_finalStep_partialProducts_T_3
    , 3'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 97:22]
  wire [4:0] quotient_finalGuess_finalStep_partialProducts_compare_4 = quotient_finalGuess_secondStep[4] ? 5'h1f : 5'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 96:24]
  wire [4:0] _quotient_finalGuess_finalStep_partialProducts_T_4 = quotient_secondGuess[4:0] &
    quotient_finalGuess_finalStep_partialProducts_compare_4; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 97:11]
  wire [8:0] quotient_finalGuess_finalStep_partialProducts_4 = {_quotient_finalGuess_finalStep_partialProducts_T_4
    , 4'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 97:22]
  wire [5:0] _GEN_27 = {{1'd0}, quotient_finalGuess_finalStep_partialProducts_0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 107:34]
  wire [6:0] _quotient_finalGuess_finalStep_partialSums_T = _GEN_27 + quotient_finalGuess_finalStep_partialProducts_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 107:34]
  wire [7:0] quotient_finalGuess_finalStep_partialSums_0 = _quotient_finalGuess_finalStep_partialSums_T +
    quotient_finalGuess_finalStep_partialProducts_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 107:39]
  wire [8:0] _GEN_28 = {{1'd0}, quotient_finalGuess_finalStep_partialProducts_3}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 108:31]
  wire [9:0] quotient_finalGuess_finalStep_partialSums_1 = _GEN_28 + quotient_finalGuess_finalStep_partialProducts_4; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 108:31]
  wire [9:0] _GEN_29 = {{2'd0}, quotient_finalGuess_finalStep_partialSums_0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:15]
  wire [10:0] _quotient_finalGuess_finalStep_T = _GEN_29 + quotient_finalGuess_finalStep_partialSums_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 104:15]
  wire [9:0] quotient_finalGuess_finalStep = _quotient_finalGuess_finalStep_T[9:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 213:27 214:17]
  wire  _quotient_finalGuess_res_roundedValue_T_4 = quotient_finalGuess_finalStep[3] & |quotient_finalGuess_finalStep[2:
    1]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 72:59]
  wire [4:0] _GEN_30 = {{4'd0}, _quotient_finalGuess_res_roundedValue_T_4}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 72:35]
  wire [5:0] quotient_finalGuess = quotient_finalGuess_finalStep[8:4] + _GEN_30; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 72:35]
  wire [2:0] dividendFraction = _shiftedValue_T[2:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 56:28 60:18]
  wire [4:0] quotient_partialProducts_compare = dividendFraction[0] ? 5'h1f : 5'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 96:24]
  wire [4:0] quotient_partialProducts_0 = quotient_finalGuess[4:0] & quotient_partialProducts_compare; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 97:11]
  wire [4:0] quotient_partialProducts_compare_1 = dividendFraction[1] ? 5'h1f : 5'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 96:24]
  wire [4:0] _quotient_partialProducts_T_1 = quotient_finalGuess[4:0] & quotient_partialProducts_compare_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 97:11]
  wire [5:0] quotient_partialProducts_1 = {_quotient_partialProducts_T_1, 1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 97:22]
  wire [4:0] quotient_partialProducts_compare_2 = dividendFraction[2] ? 5'h1f : 5'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 96:24]
  wire [4:0] _quotient_partialProducts_T_2 = quotient_finalGuess[4:0] & quotient_partialProducts_compare_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 97:11]
  wire [6:0] quotient_partialProducts_2 = {_quotient_partialProducts_T_2, 2'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 97:22]
  wire [5:0] _GEN_31 = {{1'd0}, quotient_partialProducts_0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 107:34]
  wire [6:0] _quotient_partialSums_T = _GEN_31 + quotient_partialProducts_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 107:34]
  wire [7:0] quotient = _quotient_partialSums_T + quotient_partialProducts_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 107:39]
  wire [6:0] _leadingZeros_T_39 = {quotient[0],quotient[1],quotient[2],quotient[3],quotient[4],quotient[5],quotient[6]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 58:44]
  wire [2:0] _leadingZeros_T_47 = _leadingZeros_T_39[5] ? 3'h5 : 3'h6; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] _leadingZeros_T_48 = _leadingZeros_T_39[4] ? 3'h4 : _leadingZeros_T_47; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] _leadingZeros_T_49 = _leadingZeros_T_39[3] ? 3'h3 : _leadingZeros_T_48; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] _leadingZeros_T_50 = _leadingZeros_T_39[2] ? 3'h2 : _leadingZeros_T_49; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] _leadingZeros_T_51 = _leadingZeros_T_39[1] ? 3'h1 : _leadingZeros_T_50; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] shift = _leadingZeros_T_39[0] ? 3'h0 : _leadingZeros_T_51; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [13:0] _GEN_11 = {{7'd0}, quotient[6:0]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 60:27]
  wire [13:0] _shiftedValue_T_2 = _GEN_11 << shift; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 60:27]
  wire [6:0] exponentShiftRight = 7'h0 - exponent_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 333:58]
  wire [6:0] exponentShiftLeft = exponent_1 - 7'h1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 335:38]
  wire  _T_2 = ~exponent_1[6]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 343:10]
  wire  _T_5 = ~exponent_1[6] & exponent_1[5:0] >= 6'h1f; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 343:40]
  wire  _T_12 = _T_2 & exponent_1[5:0] < 6'h1f; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 347:46]
  wire [5:0] _tempExponent_T_9 = exponent_1[5:0] + 6'h1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 349:51]
  wire [5:0] _GEN_32 = {{3'd0}, shift}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 357:78]
  wire  _T_19 = _T_2 & exponent_1[5:0] > _GEN_32; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 357:46]
  wire [6:0] shiftedCalcValue = _shiftedValue_T_2[6:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 56:28 60:18]
  wire [5:0] _tempExponent_T_12 = exponent_1[5:0] - _GEN_32; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 359:51]
  wire [132:0] _GEN_12 = {{127'd0}, quotient[6:1]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 375:83]
  wire [132:0] _tempFraction_T_3 = _GEN_12 << exponentShiftLeft; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 375:83]
  wire  _tempFraction_T_6 = &quotient[1:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 379:125]
  wire [5:0] _GEN_34 = {{5'd0}, _tempFraction_T_6}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 378:118]
  wire [5:0] _tempFraction_T_8 = quotient[7:2] + _GEN_34; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 378:118]
  wire [5:0] _tempFraction_T_9 = _tempFraction_T_8 >> exponentShiftRight; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 379:138]
  wire [132:0] _GEN_4 = _T_2 & exponent_1[5:0] > 6'h0 ? _tempFraction_T_3 : {{127'd0}, _tempFraction_T_9}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 369:82 370:22 378:22]
  wire [5:0] _GEN_5 = _T_19 & shiftedCalcValue[6] ? _tempExponent_T_12 : 6'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 358:55 359:20 368:20]
  wire [132:0] _GEN_6 = _T_19 & shiftedCalcValue[6] ? {{127'd0}, shiftedCalcValue[6:1]} : _GEN_4; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 358:55 360:20]
  wire [5:0] _GEN_7 = _T_12 & quotient[7] ? _tempExponent_T_9 : _GEN_5; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 348:54 349:20]
  wire [132:0] _GEN_8 = _T_12 & quotient[7] ? {{127'd0}, quotient[6:1]} : _GEN_6; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 348:54 350:20]
  wire [5:0] tempExponent_1 = _T_5 & quotient[7] ? 6'h1f : _GEN_7; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 344:54 345:20]
  wire [132:0] _GEN_10 = _T_5 & quotient[7] ? 133'h7f : _GEN_8; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 344:54 346:20]
  wire [6:0] tempFraction = _GEN_10[6:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 339:28]
  wire  _addOne_T_2 = roundingMode == 2'h0 & tempFraction[2]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 229:42]
  wire  _addOne_T_17 = _addOne_T_2 & ~tempFraction[1] & ~tempFraction[0] & tempFraction[3]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 230:90]
  wire  _addOne_T_18 = roundingMode == 2'h0 & tempFraction[2] & (tempFraction[1] | tempFraction[0]) | _addOne_T_17; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 229:102]
  wire  _addOne_T_24 = tempFraction[2] | tempFraction[1] | tempFraction[0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 231:70]
  wire  _addOne_T_27 = roundingMode == 2'h1 & (tempFraction[2] | tempFraction[1] | tempFraction[0]) & resultSign; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 231:90]
  wire  _addOne_T_28 = _addOne_T_18 | _addOne_T_27; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 230:110]
  wire  _addOne_T_38 = roundingMode == 2'h2 & _addOne_T_24 & ~resultSign; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 232:90]
  wire  addOne = _addOne_T_28 | _addOne_T_38; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 231:106]
  wire [2:0] _GEN_35 = {{2'd0}, addOne}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 234:66]
  wire [3:0] roundedFraction = tempFraction[5:3] + _GEN_35; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 234:66]
  wire [2:0] resultFraction = roundedFraction[3] ? roundedFraction[3:1] : roundedFraction[2:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 236:28]
  wire [5:0] _finalExponent_T_7 = tempExponent_1 + 6'h1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 240:20]
  wire [5:0] resultExponent = roundedFraction[3] | roundedFraction[2] & tempExponent_1 == 6'h0 ? _finalExponent_T_7 :
    tempExponent_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 239:28]
  wire  resultOverflow = resultExponent >= 6'h20 | tempExponent_1 == 6'h1f; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 243:59]
  assign sign = enable & resultSign; // @[\\src\\main\\scala\\fpu8\\Divide.scala 25:24 26:10 35:10]
  assign exponent = enable ? resultExponent : 6'h0; // @[\\src\\main\\scala\\fpu8\\Divide.scala 25:24 27:14 36:14]
  assign fraction = enable ? resultFraction : 3'h0; // @[\\src\\main\\scala\\fpu8\\Divide.scala 25:24 28:14 37:14]
  assign overflow = enable & resultOverflow; // @[\\src\\main\\scala\\fpu8\\Divide.scala 25:24 29:14 38:14]
  assign isInfty = enable & isResultInfty; // @[\\src\\main\\scala\\fpu8\\Divide.scala 25:24 30:13 39:13]
  assign is0 = enable & isResult0; // @[\\src\\main\\scala\\fpu8\\Divide.scala 25:24 31:9 40:9]
  assign isNaN = enable & isResultNaN; // @[\\src\\main\\scala\\fpu8\\Divide.scala 25:24 32:11 41:11]
  assign NaNFractionValue = enable & resultNaNFractionValue; // @[\\src\\main\\scala\\fpu8\\Divide.scala 25:24 33:22 42:22]
endmodule
module Compare(
  input        enable, // @[\\src\\main\\scala\\fpu8\\Compare.scala 6:18]
  input  [2:0] compareMode, // @[\\src\\main\\scala\\fpu8\\Compare.scala 7:23]
  input  [7:0] a_data, // @[\\src\\main\\scala\\fpu8\\Compare.scala 8:13]
  input  [7:0] b_data, // @[\\src\\main\\scala\\fpu8\\Compare.scala 9:13]
  output [7:0] z // @[\\src\\main\\scala\\fpu8\\Compare.scala 10:13]
);
  wire  _z_isResultNaN_T_1 = a_data[6:2] == 5'h1f; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 35:41]
  wire  _z_isResultNaN_T_3 = a_data[1:0] == 2'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 37:44]
  wire  _z_isResultNaN_T_4 = ~_z_isResultNaN_T_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 42:15]
  wire  _z_isResultNaN_T_5 = _z_isResultNaN_T_1 & _z_isResultNaN_T_4; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 41:30]
  wire  _z_isResultNaN_T_7 = b_data[6:2] == 5'h1f; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 35:41]
  wire  _z_isResultNaN_T_9 = b_data[1:0] == 2'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 37:44]
  wire  _z_isResultNaN_T_10 = ~_z_isResultNaN_T_9; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 42:15]
  wire  _z_isResultNaN_T_11 = _z_isResultNaN_T_7 & _z_isResultNaN_T_10; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 41:30]
  wire  z_isResultNaN = _z_isResultNaN_T_5 | _z_isResultNaN_T_11; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 478:34]
  wire  z_resultNaNFractionValue = a_data[1:0] > b_data[1:0] ? a_data[0] : b_data[0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 118:18]
  wire [7:0] _z_result_T = {6'h1f,1'h1,z_resultNaNFractionValue}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 483:22]
  wire  _z_T_7 = a_data[6:0] > b_data[6:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 29:77]
  wire  _z_T_11 = ~a_data[7]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 486:102]
  wire  _z_T_15 = ~_z_T_7; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 486:113]
  wire [7:0] _GEN_0 = a_data[7] > b_data[7] | a_data[7] & _z_T_7 | ~a_data[7] & ~_z_T_7 ? 8'h3c : 8'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 486:138 488:14 490:14]
  wire [7:0] z_result = z_isResultNaN ? _z_result_T : _GEN_0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 481:22 482:14]
  wire [7:0] _GEN_2 = a_data[7] < b_data[7] | a_data[7] & _z_T_15 | _z_T_11 & _z_T_7 ? 8'h3c : 8'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 507:139 509:14 511:14]
  wire [7:0] z_result_1 = z_isResultNaN ? _z_result_T : _GEN_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 502:22 503:14]
  wire [7:0] _GEN_4 = a_data == b_data ? 8'h3c : 8'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 528:42 530:14 532:14]
  wire [7:0] z_result_2 = z_isResultNaN ? _z_result_T : _GEN_4; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 523:23 524:14]
  wire [7:0] _z_result_T_26 = z_result ^ z_result_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 550:32]
  wire [7:0] z_result_3 = z_isResultNaN ? _z_result_T : _z_result_T_26; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 544:23 545:14 550:14]
  wire [7:0] _z_result_T_47 = z_result_1 ^ z_result_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 568:32]
  wire [7:0] z_result_4 = z_isResultNaN ? _z_result_T : _z_result_T_47; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 562:23 563:14 568:14]
  wire [7:0] _GEN_16 = a_data != b_data ? 8'h3c : 8'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 585:42 587:14 589:14]
  wire [7:0] z_result_5 = z_isResultNaN ? _z_result_T : _GEN_16; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 580:23 581:14]
  wire [7:0] _GEN_18 = compareMode == 3'h4 ? z_result_4 : z_result_5; // @[\\src\\main\\scala\\fpu8\\Compare.scala 21:37 22:9 24:9]
  wire [7:0] _GEN_19 = compareMode == 3'h3 ? z_result_3 : _GEN_18; // @[\\src\\main\\scala\\fpu8\\Compare.scala 19:37 20:9]
  wire [7:0] _GEN_20 = compareMode == 3'h2 ? z_result_2 : _GEN_19; // @[\\src\\main\\scala\\fpu8\\Compare.scala 17:37 18:9]
  wire [7:0] _GEN_21 = compareMode == 3'h1 ? z_result_1 : _GEN_20; // @[\\src\\main\\scala\\fpu8\\Compare.scala 15:37 16:9]
  wire [7:0] _GEN_22 = compareMode == 3'h0 ? z_result : _GEN_21; // @[\\src\\main\\scala\\fpu8\\Compare.scala 13:31 14:9]
  assign z = enable ? _GEN_22 : 8'h0; // @[\\src\\main\\scala\\fpu8\\Compare.scala 12:23 27:6]
endmodule
module Convert(
  input        enable, // @[\\src\\main\\scala\\fpu8\\Convert.scala 6:18]
  input  [7:0] a_data, // @[\\src\\main\\scala\\fpu8\\Convert.scala 7:13]
  input  [1:0] roundingMode, // @[\\src\\main\\scala\\fpu8\\Convert.scala 8:24]
  input        saturationMode, // @[\\src\\main\\scala\\fpu8\\Convert.scala 9:26]
  output [7:0] z // @[\\src\\main\\scala\\fpu8\\Convert.scala 10:13]
);
  wire  _z_isResultNaN_T_1 = a_data[6:2] == 5'h1f; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 35:41]
  wire  _z_isResultNaN_T_3 = a_data[1:0] == 2'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 37:44]
  wire  _z_isResultNaN_T_4 = ~_z_isResultNaN_T_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 42:15]
  wire  _z_isResultNaN_T_5 = _z_isResultNaN_T_1 & _z_isResultNaN_T_4; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 41:30]
  wire  _z_isResultNaN_T_10 = _z_isResultNaN_T_1 & _z_isResultNaN_T_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 47:24]
  wire  z_isResultNaN = _z_isResultNaN_T_5 | _z_isResultNaN_T_10; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 628:29]
  wire  _z_fraction_T_1 = a_data[6:2] == 5'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 33:39]
  wire  _z_fraction_T_2 = ~_z_fraction_T_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 630:24]
  wire [5:0] z_tempExponent = a_data[6:2] - 5'h8; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 632:33]
  wire  z_isDenormalized = z_tempExponent[5] | z_tempExponent[4:0] == 5'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 634:55]
  wire  z_overflow = ~z_tempExponent[5] & z_tempExponent[4]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 635:50]
  wire [6:0] _z_shift_T = 6'h1 - z_tempExponent; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 636:41]
  wire [6:0] z_shift = z_isDenormalized ? _z_shift_T : 7'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 636:20]
  wire [6:0] _z_tempFraction_T = {_z_fraction_T_2,a_data[1:0],4'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 638:27]
  wire [6:0] z_tempFraction = _z_tempFraction_T >> z_shift; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 638:67]
  wire  _z_addOne_T = roundingMode == 2'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 640:33]
  wire  _z_addOne_T_2 = roundingMode == 2'h0 & z_tempFraction[2]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 640:42]
  wire  _z_addOne_T_17 = _z_addOne_T_2 & ~z_tempFraction[1] & ~z_tempFraction[0] & z_tempFraction[3]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 641:90]
  wire  _z_addOne_T_18 = roundingMode == 2'h0 & z_tempFraction[2] & (z_tempFraction[1] | z_tempFraction[0]) |
    _z_addOne_T_17; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 640:102]
  wire  _z_addOne_T_19 = roundingMode == 2'h1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 642:22]
  wire  _z_addOne_T_24 = z_tempFraction[2] | z_tempFraction[1] | z_tempFraction[0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 642:70]
  wire  _z_addOne_T_28 = roundingMode == 2'h1 & (z_tempFraction[2] | z_tempFraction[1] | z_tempFraction[0]) & a_data[7]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 642:90]
  wire  _z_addOne_T_29 = _z_addOne_T_18 | _z_addOne_T_28; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 641:110]
  wire  _z_addOne_T_30 = roundingMode == 2'h2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 643:22]
  wire  _z_addOne_T_39 = ~a_data[7]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 643:93]
  wire  _z_addOne_T_40 = roundingMode == 2'h2 & _z_addOne_T_24 & ~a_data[7]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 643:90]
  wire  z_addOne = _z_addOne_T_29 | _z_addOne_T_40; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 642:106]
  wire [3:0] _GEN_8 = {{3'd0}, z_addOne}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 645:80]
  wire [4:0] z_roundedFraction = z_tempFraction[6:3] + _GEN_8; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 645:80]
  wire [3:0] _z_finalExponent_T_1 = z_isDenormalized ? 4'h0 : z_tempExponent[3:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 648:10]
  wire [3:0] z_finalExponent = z_overflow ? 4'hf : _z_finalExponent_T_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 647:28]
  wire [3:0] z_finalFraction = z_roundedFraction[3:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 650:40]
  wire  _z_T_2 = ~saturationMode; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 656:54]
  wire  _z_T_9 = _z_addOne_T_19 & _z_T_2 & _z_addOne_T_39; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 657:59]
  wire  _z_T_10 = _z_addOne_T & ~saturationMode | _z_T_9; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 656:63]
  wire  _z_T_16 = _z_addOne_T_30 & _z_T_2 & _z_addOne_T_39; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 658:59]
  wire  _z_T_17 = _z_T_10 | _z_T_16; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 657:76]
  wire  _z_T_23 = roundingMode == 2'h3 & _z_T_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 661:33]
  wire  _z_T_24 = _z_addOne_T & saturationMode | _z_T_23; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 660:69]
  wire [7:0] _z_result_T_2 = {a_data[7],4'hf,3'h6}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 662:24]
  wire  _z_T_34 = _z_addOne_T_30 & a_data[7]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 664:33]
  wire  _z_T_35 = _z_addOne_T_19 & saturationMode & _z_addOne_T_39 | _z_T_34; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 663:85]
  wire  _z_T_45 = _z_addOne_T_30 & saturationMode & _z_addOne_T_39; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 667:59]
  wire  _z_T_46 = _z_addOne_T_19 & a_data[7] | _z_T_45; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 666:59]
  wire [7:0] _GEN_0 = _z_T_46 ? _z_result_T_2 : 8'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 667:77 668:18 670:18]
  wire [7:0] _GEN_1 = _z_T_35 ? _z_result_T_2 : _GEN_0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 664:51 665:18]
  wire [7:0] _GEN_2 = _z_T_24 ? _z_result_T_2 : _GEN_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 661:61 662:18]
  wire [7:0] _GEN_3 = _z_T_17 ? 8'h7f : _GEN_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 658:77 659:18]
  wire [7:0] _z_result_T_9 = {a_data[7],z_finalExponent,z_finalFraction[2:0]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 673:22]
  wire [7:0] _GEN_4 = z_overflow ? _GEN_3 : _z_result_T_9; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 655:22 673:16]
  wire [7:0] _GEN_5 = z_isResultNaN ? 8'h7f : 8'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 675:29 676:14 678:14]
  wire [7:0] z_result = ~z_isResultNaN ? _GEN_4 : _GEN_5; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 654:24]
  assign z = enable ? z_result : 8'h0; // @[\\src\\main\\scala\\fpu8\\Convert.scala 12:23 13:7 18:7]
endmodule
module GenerateFinalResult(
  input        enable, // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 12:18]
  input        sign, // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 13:16]
  input  [4:0] exponent, // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 14:20]
  input  [1:0] mantissa, // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 15:20]
  input  [1:0] roundingMode, // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 16:24]
  input        overflow, // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 17:20]
  input        saturationMode, // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 18:26]
  input        isInfty, // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 19:19]
  input        is0, // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 20:15]
  input        isNaN, // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 21:17]
  input        NaNFractionValue, // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 22:28]
  output [7:0] z // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 23:13]
);
  wire  _result_T_4 = ~isInfty; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 70:10]
  wire  _result_T_5 = ~is0; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 70:22]
  wire  _result_T_7 = ~isNaN; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 70:30]
  wire  _result_T_9 = roundingMode == 2'h0; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 72:27]
  wire  _result_T_10 = ~saturationMode; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 72:53]
  wire [7:0] _result_z_T = {sign,5'h1f,2'h0}; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 73:19]
  wire [7:0] _result_z_T_1 = {sign,5'h1e,2'h3}; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 75:19]
  wire  _result_T_17 = roundingMode == 2'h1; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 76:33]
  wire  _result_T_20 = ~sign; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 76:75]
  wire  _result_T_27 = roundingMode == 2'h2; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 78:102]
  wire [7:0] _GEN_0 = _result_T_27 & _result_T_10 & _result_T_20 ? 8'h7c : 8'h0; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 82:84 83:13 85:13]
  wire [7:0] _GEN_1 = _result_T_17 & sign | _result_T_27 & saturationMode & _result_T_20 ? 8'h7b : _GEN_0; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 80:128 81:13]
  wire [7:0] _GEN_2 = _result_T_17 & saturationMode & _result_T_20 | roundingMode == 2'h2 & sign ? 8'hfb : _GEN_1; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 78:128 79:13]
  wire [7:0] _GEN_3 = roundingMode == 2'h1 & _result_T_10 & ~sign ? 8'hfc : _GEN_2; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 76:84 77:13]
  wire [7:0] _GEN_4 = _result_T_9 & saturationMode | roundingMode == 2'h3 ? _result_z_T_1 : _GEN_3; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 74:94 75:13]
  wire [7:0] _GEN_5 = roundingMode == 2'h0 & ~saturationMode ? _result_z_T : _GEN_4; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 72:62 73:13]
  wire [7:0] _result_z_T_6 = {sign,exponent,mantissa}; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 88:17]
  wire [7:0] _GEN_6 = overflow ? _GEN_5 : _result_z_T_6; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 71:22 88:11]
  wire [7:0] _result_z_T_8 = {sign,5'h0,2'h0}; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 93:15]
  wire [7:0] _result_z_T_9 = {6'h1f,1'h1,NaNFractionValue}; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 95:15]
  wire [7:0] _GEN_7 = isNaN ? _result_z_T_9 : 8'h0; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 94:23 95:9 97:9]
  wire [7:0] _GEN_8 = _result_T_4 & is0 & _result_T_7 ? _result_z_T_8 : _GEN_7; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 92:43 93:9]
  wire [7:0] _GEN_9 = isInfty & _result_T_5 & _result_T_7 ? _result_z_T : _GEN_8; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 90:43 91:9]
  wire [7:0] result = ~isInfty & ~is0 & ~isNaN ? _GEN_6 : _GEN_9; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 70:38]
  assign z = enable ? result : 8'h0; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 31:23 32:7 34:7]
endmodule
module FPU8Generator(
  input        clock,
  input        reset,
  input        enable, // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 9:18]
  input  [7:0] a_data, // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 10:13]
  input  [7:0] b_data, // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 11:13]
  input  [3:0] opCode, // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 12:18]
  input  [1:0] roundingMode, // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 13:24]
  input        saturationMode, // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 14:26]
  output [7:0] z // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 15:13]
);
  wire  addSub_enable; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 17:22]
  wire [7:0] addSub_a_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 17:22]
  wire [7:0] addSub_b_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 17:22]
  wire  addSub_subtract; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 17:22]
  wire [1:0] addSub_roundingMode; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 17:22]
  wire  addSub_sign; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 17:22]
  wire [5:0] addSub_exponent; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 17:22]
  wire [2:0] addSub_fraction; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 17:22]
  wire  addSub_overflow; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 17:22]
  wire  addSub_isInfty; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 17:22]
  wire  addSub_is0; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 17:22]
  wire  addSub_isNaN; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 17:22]
  wire  addSub_NaNFractionValue; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 17:22]
  wire  multiply_enable; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 19:24]
  wire [7:0] multiply_a_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 19:24]
  wire [7:0] multiply_b_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 19:24]
  wire [1:0] multiply_roundingMode; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 19:24]
  wire  multiply_sign; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 19:24]
  wire [5:0] multiply_exponent; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 19:24]
  wire [2:0] multiply_fraction; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 19:24]
  wire  multiply_overflow; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 19:24]
  wire  multiply_isInfty; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 19:24]
  wire  multiply_is0; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 19:24]
  wire  multiply_isNaN; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 19:24]
  wire  multiply_NaNFractionValue; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 19:24]
  wire  divide_enable; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 21:22]
  wire [7:0] divide_a_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 21:22]
  wire [7:0] divide_b_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 21:22]
  wire [1:0] divide_roundingMode; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 21:22]
  wire  divide_sign; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 21:22]
  wire [5:0] divide_exponent; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 21:22]
  wire [2:0] divide_fraction; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 21:22]
  wire  divide_overflow; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 21:22]
  wire  divide_isInfty; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 21:22]
  wire  divide_is0; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 21:22]
  wire  divide_isNaN; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 21:22]
  wire  divide_NaNFractionValue; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 21:22]
  wire  compare_enable; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 23:23]
  wire [2:0] compare_compareMode; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 23:23]
  wire [7:0] compare_a_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 23:23]
  wire [7:0] compare_b_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 23:23]
  wire [7:0] compare_z; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 23:23]
  wire  convert_enable; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 25:23]
  wire [7:0] convert_a_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 25:23]
  wire [1:0] convert_roundingMode; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 25:23]
  wire  convert_saturationMode; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 25:23]
  wire [7:0] convert_z; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 25:23]
  wire  generateFinalResult_enable; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 27:35]
  wire  generateFinalResult_sign; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 27:35]
  wire [4:0] generateFinalResult_exponent; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 27:35]
  wire [1:0] generateFinalResult_mantissa; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 27:35]
  wire [1:0] generateFinalResult_roundingMode; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 27:35]
  wire  generateFinalResult_overflow; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 27:35]
  wire  generateFinalResult_saturationMode; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 27:35]
  wire  generateFinalResult_isInfty; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 27:35]
  wire  generateFinalResult_is0; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 27:35]
  wire  generateFinalResult_isNaN; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 27:35]
  wire  generateFinalResult_NaNFractionValue; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 27:35]
  wire [7:0] generateFinalResult_z; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 27:35]
  wire  _addSub_enable_T_2 = opCode == 4'h0 | opCode == 4'h1; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 29:39]
  wire  _multiply_enable_T = opCode == 4'h2; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 35:33]
  wire  _divide_enable_T = opCode == 4'h3; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 40:31]
  wire  _compare_enable_T = opCode == 4'h4; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 45:32]
  wire  _compare_enable_T_1 = opCode == 4'h5; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 45:50]
  wire  _compare_enable_T_3 = opCode == 4'h6; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 45:68]
  wire  _compare_enable_T_5 = opCode == 4'h7; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 45:86]
  wire  _compare_enable_T_7 = opCode == 4'h8; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 45:104]
  wire  _compare_enable_T_10 = opCode == 4'h4 | opCode == 4'h5 | opCode == 4'h6 | opCode == 4'h7 | opCode == 4'h8 |
    opCode == 4'h9; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 45:112]
  wire [2:0] _compare_compareMode_T_5 = _compare_enable_T_7 ? 3'h4 : 3'h5; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 51:14]
  wire [2:0] _compare_compareMode_T_6 = _compare_enable_T_5 ? 3'h3 : _compare_compareMode_T_5; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 50:12]
  wire [2:0] _compare_compareMode_T_7 = _compare_enable_T_3 ? 3'h2 : _compare_compareMode_T_6; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 49:10]
  wire [2:0] _compare_compareMode_T_8 = _compare_enable_T_1 ? 3'h1 : _compare_compareMode_T_7; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 48:8]
  wire  _convert_enable_T = opCode == 4'ha; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 55:32]
  wire [7:0] _GEN_1 = _convert_enable_T ? convert_z : 8'h0; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 114:30 126:7 139:7]
  wire [7:0] _GEN_3 = _compare_enable_T_10 ? compare_z : _GEN_1; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 101:119 113:7]
  wire  _GEN_4 = _divide_enable_T & divide_sign; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 88:30 89:30]
  wire [4:0] _GEN_5 = _divide_enable_T ? divide_exponent[4:0] : 5'h0; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 88:30 90:34]
  wire [1:0] _GEN_6 = _divide_enable_T ? divide_fraction[1:0] : 2'h0; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 88:30 91:34]
  wire [1:0] _GEN_7 = _divide_enable_T ? roundingMode : 2'h0; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 88:30 92:38]
  wire  _GEN_8 = _divide_enable_T & divide_overflow; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 88:30 93:34]
  wire  _GEN_9 = _divide_enable_T & saturationMode; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 88:30 94:40]
  wire  _GEN_10 = _divide_enable_T & divide_isInfty; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 88:30 95:33]
  wire  _GEN_11 = _divide_enable_T & divide_is0; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 88:30 96:29]
  wire  _GEN_12 = _divide_enable_T & divide_isNaN; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 88:30 97:31]
  wire  _GEN_13 = _divide_enable_T & divide_NaNFractionValue; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 88:30 98:42]
  wire [7:0] _GEN_14 = _divide_enable_T ? generateFinalResult_z : _GEN_3; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 88:30 100:7]
  wire  _GEN_15 = _multiply_enable_T ? multiply_sign : _GEN_4; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 75:30 76:30]
  wire [4:0] _GEN_16 = _multiply_enable_T ? multiply_exponent[4:0] : _GEN_5; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 75:30 77:34]
  wire [1:0] _GEN_17 = _multiply_enable_T ? multiply_fraction[1:0] : _GEN_6; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 75:30 78:34]
  wire [1:0] _GEN_18 = _multiply_enable_T ? roundingMode : _GEN_7; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 75:30 79:38]
  wire  _GEN_19 = _multiply_enable_T ? multiply_overflow : _GEN_8; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 75:30 80:34]
  wire  _GEN_20 = _multiply_enable_T ? saturationMode : _GEN_9; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 75:30 81:40]
  wire  _GEN_21 = _multiply_enable_T ? multiply_isInfty : _GEN_10; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 75:30 82:33]
  wire  _GEN_22 = _multiply_enable_T ? multiply_is0 : _GEN_11; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 75:30 83:29]
  wire  _GEN_23 = _multiply_enable_T ? multiply_isNaN : _GEN_12; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 75:30 84:31]
  wire  _GEN_24 = _multiply_enable_T ? multiply_NaNFractionValue : _GEN_13; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 75:30 85:42]
  wire [7:0] _GEN_25 = _multiply_enable_T ? generateFinalResult_z : _GEN_14; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 75:30 87:7]
  Add addSub ( // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 17:22]
    .enable(addSub_enable),
    .a_data(addSub_a_data),
    .b_data(addSub_b_data),
    .subtract(addSub_subtract),
    .roundingMode(addSub_roundingMode),
    .sign(addSub_sign),
    .exponent(addSub_exponent),
    .fraction(addSub_fraction),
    .overflow(addSub_overflow),
    .isInfty(addSub_isInfty),
    .is0(addSub_is0),
    .isNaN(addSub_isNaN),
    .NaNFractionValue(addSub_NaNFractionValue)
  );
  Multiply multiply ( // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 19:24]
    .enable(multiply_enable),
    .a_data(multiply_a_data),
    .b_data(multiply_b_data),
    .roundingMode(multiply_roundingMode),
    .sign(multiply_sign),
    .exponent(multiply_exponent),
    .fraction(multiply_fraction),
    .overflow(multiply_overflow),
    .isInfty(multiply_isInfty),
    .is0(multiply_is0),
    .isNaN(multiply_isNaN),
    .NaNFractionValue(multiply_NaNFractionValue)
  );
  Divide divide ( // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 21:22]
    .enable(divide_enable),
    .a_data(divide_a_data),
    .b_data(divide_b_data),
    .roundingMode(divide_roundingMode),
    .sign(divide_sign),
    .exponent(divide_exponent),
    .fraction(divide_fraction),
    .overflow(divide_overflow),
    .isInfty(divide_isInfty),
    .is0(divide_is0),
    .isNaN(divide_isNaN),
    .NaNFractionValue(divide_NaNFractionValue)
  );
  Compare compare ( // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 23:23]
    .enable(compare_enable),
    .compareMode(compare_compareMode),
    .a_data(compare_a_data),
    .b_data(compare_b_data),
    .z(compare_z)
  );
  Convert convert ( // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 25:23]
    .enable(convert_enable),
    .a_data(convert_a_data),
    .roundingMode(convert_roundingMode),
    .saturationMode(convert_saturationMode),
    .z(convert_z)
  );
  GenerateFinalResult generateFinalResult ( // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 27:35]
    .enable(generateFinalResult_enable),
    .sign(generateFinalResult_sign),
    .exponent(generateFinalResult_exponent),
    .mantissa(generateFinalResult_mantissa),
    .roundingMode(generateFinalResult_roundingMode),
    .overflow(generateFinalResult_overflow),
    .saturationMode(generateFinalResult_saturationMode),
    .isInfty(generateFinalResult_isInfty),
    .is0(generateFinalResult_is0),
    .isNaN(generateFinalResult_isNaN),
    .NaNFractionValue(generateFinalResult_NaNFractionValue),
    .z(generateFinalResult_z)
  );
  assign z = _addSub_enable_T_2 ? generateFinalResult_z : _GEN_25; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 62:42 74:7]
  assign addSub_enable = (opCode == 4'h0 | opCode == 4'h1) & enable; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 29:23]
  assign addSub_a_data = a_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 30:12]
  assign addSub_b_data = b_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 31:12]
  assign addSub_subtract = opCode == 4'h1; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 32:33]
  assign addSub_roundingMode = roundingMode; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 33:23]
  assign multiply_enable = opCode == 4'h2 & enable; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 35:25]
  assign multiply_a_data = a_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 36:14]
  assign multiply_b_data = b_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 37:14]
  assign multiply_roundingMode = roundingMode; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 38:25]
  assign divide_enable = opCode == 4'h3 & enable; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 40:23]
  assign divide_a_data = a_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 41:12]
  assign divide_b_data = b_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 42:12]
  assign divide_roundingMode = roundingMode; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 43:23]
  assign compare_enable = (opCode == 4'h4 | opCode == 4'h5 | opCode == 4'h6 | opCode == 4'h7 | opCode == 4'h8 | opCode
     == 4'h9) & enable; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 45:24]
  assign compare_compareMode = _compare_enable_T ? 3'h0 : _compare_compareMode_T_8; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 47:29]
  assign compare_a_data = a_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 52:13]
  assign compare_b_data = b_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 53:13]
  assign convert_enable = opCode == 4'ha & enable; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 55:24]
  assign convert_a_data = a_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 56:13]
  assign convert_roundingMode = roundingMode; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 57:24]
  assign convert_saturationMode = saturationMode; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 58:26]
  assign generateFinalResult_enable = enable; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 60:30]
  assign generateFinalResult_sign = _addSub_enable_T_2 ? addSub_sign : _GEN_15; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 62:42 63:30]
  assign generateFinalResult_exponent = _addSub_enable_T_2 ? addSub_exponent[4:0] : _GEN_16; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 62:42 64:34]
  assign generateFinalResult_mantissa = _addSub_enable_T_2 ? addSub_fraction[1:0] : _GEN_17; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 62:42 65:34]
  assign generateFinalResult_roundingMode = _addSub_enable_T_2 ? roundingMode : _GEN_18; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 62:42 66:38]
  assign generateFinalResult_overflow = _addSub_enable_T_2 ? addSub_overflow : _GEN_19; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 62:42 67:34]
  assign generateFinalResult_saturationMode = _addSub_enable_T_2 ? saturationMode : _GEN_20; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 62:42 68:40]
  assign generateFinalResult_isInfty = _addSub_enable_T_2 ? addSub_isInfty : _GEN_21; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 62:42 69:33]
  assign generateFinalResult_is0 = _addSub_enable_T_2 ? addSub_is0 : _GEN_22; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 62:42 70:29]
  assign generateFinalResult_isNaN = _addSub_enable_T_2 ? addSub_isNaN : _GEN_23; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 62:42 71:31]
  assign generateFinalResult_NaNFractionValue = _addSub_enable_T_2 ? addSub_NaNFractionValue : _GEN_24; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 62:42 72:42]
endmodule
