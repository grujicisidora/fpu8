module Add(
  input        enable, // @[\\src\\main\\scala\\fpu8\\Add.scala 10:18]
  input  [7:0] a_data, // @[\\src\\main\\scala\\fpu8\\Add.scala 11:13]
  input  [7:0] b_data, // @[\\src\\main\\scala\\fpu8\\Add.scala 12:13]
  input        subtract, // @[\\src\\main\\scala\\fpu8\\Add.scala 13:20]
  input  [1:0] roundingMode, // @[\\src\\main\\scala\\fpu8\\Add.scala 14:24]
  output       sign, // @[\\src\\main\\scala\\fpu8\\Add.scala 15:16]
  output [5:0] exponent, // @[\\src\\main\\scala\\fpu8\\Add.scala 16:20]
  output [2:0] fraction, // @[\\src\\main\\scala\\fpu8\\Add.scala 17:20]
  output       NaNFractionValue, // @[\\src\\main\\scala\\fpu8\\Add.scala 18:28]
  output [4:0] status // @[\\src\\main\\scala\\fpu8\\Add.scala 19:18]
);
  wire  compare = a_data[6:0] > b_data[6:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 29:77]
  wire [7:0] greaterOperand_data = compare ? a_data : b_data; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 129:29]
  wire [7:0] smallerOperand_data = compare ? b_data : a_data; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 130:29]
  wire  resultSign = compare ? a_data[7] : b_data[7] ^ subtract; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 131:19]
  wire  subtraction = subtract ^ greaterOperand_data[7] ^ smallerOperand_data[7]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 132:54]
  wire [4:0] exponent_1 = greaterOperand_data[6:2]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 25:28]
  wire  _greaterOperandFraction_T_1 = exponent_1 == 5'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 33:39]
  wire  _greaterOperandFraction_T_2 = ~_greaterOperandFraction_T_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 134:38]
  wire  _smallerOperandFraction_T_1 = smallerOperand_data[6:2] == 5'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 33:39]
  wire  _smallerOperandFraction_T_2 = ~_smallerOperandFraction_T_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 135:38]
  wire  isOnlySmallerDenormalized = _greaterOperandFraction_T_2 & _smallerOperandFraction_T_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 136:60]
  wire [4:0] _shift_T_2 = exponent_1 - 5'h1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 139:31]
  wire [4:0] _shift_T_6 = exponent_1 - smallerOperand_data[6:2]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 140:31]
  wire [4:0] shift = isOnlySmallerDenormalized ? _shift_T_2 : _shift_T_6; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 137:20]
  wire  _shiftedFraction_shifted_T = shift >= 5'h5; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 145:15]
  wire [7:0] _shiftedFraction_shifted_T_1 = {5'h0,_smallerOperandFraction_T_2,smallerOperand_data[1:0]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 146:12]
  wire [7:0] _shiftedFraction_shifted_T_2 = {_smallerOperandFraction_T_2,smallerOperand_data[1:0],5'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 147:12]
  wire [7:0] _shiftedFraction_shifted_T_3 = _shiftedFraction_shifted_T_2 >> shift; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 147:54]
  wire [7:0] shiftedFraction_shifted = _shiftedFraction_shifted_T ? _shiftedFraction_shifted_T_1 :
    _shiftedFraction_shifted_T_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 144:24]
  wire [5:0] smallerOperandFraction_1 = {shiftedFraction_shifted[7:3],|shiftedFraction_shifted[2:0]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 149:10]
  wire [5:0] greaterOperandFraction_1 = {_greaterOperandFraction_T_2,greaterOperand_data[1:0],3'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 151:45]
  wire  _isResultNaN_T_1 = a_data[6:2] == 5'h1f; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 35:41]
  wire  _isResultNaN_T_3 = a_data[1:0] == 2'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 37:44]
  wire  _isResultNaN_T_4 = ~_isResultNaN_T_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 42:15]
  wire  _isResultNaN_T_5 = _isResultNaN_T_1 & _isResultNaN_T_4; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 41:30]
  wire  _isResultNaN_T_7 = b_data[6:2] == 5'h1f; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 35:41]
  wire  _isResultNaN_T_9 = b_data[1:0] == 2'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 37:44]
  wire  _isResultNaN_T_10 = ~_isResultNaN_T_9; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 42:15]
  wire  _isResultNaN_T_11 = _isResultNaN_T_7 & _isResultNaN_T_10; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 41:30]
  wire  _isResultNaN_T_17 = _isResultNaN_T_1 & _isResultNaN_T_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 47:24]
  wire  _isResultNaN_T_22 = _isResultNaN_T_7 & _isResultNaN_T_9; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 47:24]
  wire  isResultNaN = _isResultNaN_T_5 | _isResultNaN_T_11 | _isResultNaN_T_17 & _isResultNaN_T_22 & subtraction; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 413:57]
  wire  _isResultInfty_T_11 = ~isResultNaN; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 418:65]
  wire  isResultInfty = (_isResultNaN_T_17 | _isResultNaN_T_22) & ~isResultNaN; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 418:63]
  wire  _isResult0_T_2 = a_data[6:0] == b_data[6:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 31:77]
  wire  isResult0 = _isResult0_T_2 & subtraction & _isResultInfty_T_11 & ~isResultInfty; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 422:101]
  wire  resultNaNFractionValue = a_data[1:0] > b_data[1:0] ? a_data[0] : b_data[0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 123:18]
  wire [6:0] _calculatedValue_T_1 = greaterOperandFraction_1 - smallerOperandFraction_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 427:32]
  wire [6:0] _calculatedValue_T_3 = greaterOperandFraction_1 + smallerOperandFraction_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 428:32]
  wire [6:0] calculatedValue = subtraction ? _calculatedValue_T_1 : _calculatedValue_T_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 426:32]
  wire [7:0] paddedCalcValue = {calculatedValue,1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 267:15]
  wire [6:0] _leadingZeros_T_17 = {paddedCalcValue[0],paddedCalcValue[1],paddedCalcValue[2],paddedCalcValue[3],
    paddedCalcValue[4],paddedCalcValue[5],paddedCalcValue[6]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 58:44]
  wire [2:0] _leadingZeros_T_25 = _leadingZeros_T_17[5] ? 3'h5 : 3'h6; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] _leadingZeros_T_26 = _leadingZeros_T_17[4] ? 3'h4 : _leadingZeros_T_25; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] _leadingZeros_T_27 = _leadingZeros_T_17[3] ? 3'h3 : _leadingZeros_T_26; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] _leadingZeros_T_28 = _leadingZeros_T_17[2] ? 3'h2 : _leadingZeros_T_27; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] _leadingZeros_T_29 = _leadingZeros_T_17[1] ? 3'h1 : _leadingZeros_T_28; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] shift_1 = _leadingZeros_T_17[0] ? 3'h0 : _leadingZeros_T_29; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [7:0] _shiftedValue_T_3 = {paddedCalcValue[6:0], 1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 63:23]
  wire [8:0] _shiftedValue_T_5 = {paddedCalcValue[6:0], 2'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 63:23]
  wire [9:0] _shiftedValue_T_7 = {paddedCalcValue[6:0], 3'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 63:23]
  wire [10:0] _shiftedValue_T_9 = {paddedCalcValue[6:0], 4'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 63:23]
  wire [11:0] _shiftedValue_T_11 = {paddedCalcValue[6:0], 5'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 63:23]
  wire [12:0] _shiftedValue_T_13 = {paddedCalcValue[6:0], 6'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 63:23]
  wire [6:0] _shiftedValue_T_18 = 3'h1 == shift_1 ? _shiftedValue_T_3[6:0] : paddedCalcValue[6:0]; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [6:0] _shiftedValue_T_20 = 3'h2 == shift_1 ? _shiftedValue_T_5[6:0] : _shiftedValue_T_18; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [6:0] _shiftedValue_T_22 = 3'h3 == shift_1 ? _shiftedValue_T_7[6:0] : _shiftedValue_T_20; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [6:0] _shiftedValue_T_24 = 3'h4 == shift_1 ? _shiftedValue_T_9[6:0] : _shiftedValue_T_22; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [6:0] _shiftedValue_T_26 = 3'h5 == shift_1 ? _shiftedValue_T_11[6:0] : _shiftedValue_T_24; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [6:0] shiftedCalcValue = 3'h6 == shift_1 ? _shiftedValue_T_13[6:0] : _shiftedValue_T_26; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire  _T_1 = &exponent_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 275:19]
  wire [4:0] _tempExponent_T_1 = exponent_1 + 5'h1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 279:32]
  wire [6:0] _tempFraction_T_3 = {paddedCalcValue[7:2],|paddedCalcValue[1:0]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 280:26]
  wire [4:0] _GEN_12 = {{2'd0}, shift_1}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 281:25]
  wire [4:0] _tempExponent_T_3 = exponent_1 - _GEN_12; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 282:32]
  wire [37:0] _GEN_5 = {{31'd0}, paddedCalcValue[6:0]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 287:47]
  wire [37:0] _tempFraction_T_7 = _GEN_5 << _shift_T_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 287:47]
  wire [37:0] _GEN_0 = exponent_1 > 5'h0 ? _tempFraction_T_7 : {{31'd0}, paddedCalcValue[6:0]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 286:28 287:22 289:22]
  wire [4:0] _GEN_1 = exponent_1 > _GEN_12 & shiftedCalcValue[6] ? _tempExponent_T_3 : 5'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 281:57 282:20 285:20]
  wire [37:0] _GEN_2 = exponent_1 > _GEN_12 & shiftedCalcValue[6] ? {{31'd0}, shiftedCalcValue} : _GEN_0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 281:57 283:20]
  wire [4:0] _GEN_3 = ~_T_1 & paddedCalcValue[7] ? _tempExponent_T_1 : _GEN_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 278:54 279:20]
  wire [37:0] _GEN_4 = ~_T_1 & paddedCalcValue[7] ? {{31'd0}, _tempFraction_T_3} : _GEN_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 278:54 280:20]
  wire [4:0] tempExponent = &exponent_1 & paddedCalcValue[7] ? exponent_1 : _GEN_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 275:47 276:20]
  wire [37:0] _GEN_6 = &exponent_1 & paddedCalcValue[7] ? 38'h7f : _GEN_4; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 275:47 277:20]
  wire [6:0] tempFraction = _GEN_6[6:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 273:28]
  wire  _addOne_T_2 = roundingMode == 2'h0 & tempFraction[3]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 234:42]
  wire  _addOne_T_17 = _addOne_T_2 & ~tempFraction[2] & ~tempFraction[1] & tempFraction[4]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 235:90]
  wire  _addOne_T_18 = roundingMode == 2'h0 & tempFraction[3] & (tempFraction[2] | tempFraction[1]) | _addOne_T_17; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 234:102]
  wire  _addOne_T_24 = tempFraction[3] | tempFraction[2] | tempFraction[1]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 236:70]
  wire  _addOne_T_27 = roundingMode == 2'h1 & (tempFraction[3] | tempFraction[2] | tempFraction[1]) & resultSign; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 236:90]
  wire  _addOne_T_28 = _addOne_T_18 | _addOne_T_27; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 235:110]
  wire  _addOne_T_38 = roundingMode == 2'h2 & _addOne_T_24 & ~resultSign; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 237:90]
  wire  addOne = _addOne_T_28 | _addOne_T_38; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 236:106]
  wire [2:0] _GEN_14 = {{2'd0}, addOne}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 239:66]
  wire [3:0] roundedFraction = tempFraction[6:4] + _GEN_14; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 239:66]
  wire [2:0] resultFraction = roundedFraction[3] ? roundedFraction[3:1] : roundedFraction[2:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 241:28]
  wire [4:0] _finalExponent_T_7 = tempExponent + 5'h1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 245:20]
  wire [4:0] resultExponent = roundedFraction[3] | roundedFraction[2] & tempExponent == 5'h0 ? _finalExponent_T_7 :
    tempExponent; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 244:28]
  wire  overflow = tempExponent == 5'h1f; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 248:76]
  wire [4:0] resultStatus = {overflow,resultExponent == 5'h0,isResultNaN,isResultInfty,isResult0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 432:23]
  wire [4:0] _GEN_8 = enable ? resultExponent : 5'h0; // @[\\src\\main\\scala\\fpu8\\Add.scala 24:24 26:14 32:14]
  assign sign = enable & resultSign; // @[\\src\\main\\scala\\fpu8\\Add.scala 24:24 25:10 31:10]
  assign exponent = {{1'd0}, _GEN_8};
  assign fraction = enable ? resultFraction : 3'h0; // @[\\src\\main\\scala\\fpu8\\Add.scala 24:24 27:14 33:14]
  assign NaNFractionValue = enable & resultNaNFractionValue; // @[\\src\\main\\scala\\fpu8\\Add.scala 24:24 29:22 35:22]
  assign status = enable ? resultStatus : 5'h0; // @[\\src\\main\\scala\\fpu8\\Add.scala 24:24 28:12 34:12]
endmodule
module Multiply(
  input        enable, // @[\\src\\main\\scala\\fpu8\\Multiply.scala 10:18]
  input  [7:0] a_data, // @[\\src\\main\\scala\\fpu8\\Multiply.scala 11:13]
  input  [7:0] b_data, // @[\\src\\main\\scala\\fpu8\\Multiply.scala 12:13]
  input  [1:0] roundingMode, // @[\\src\\main\\scala\\fpu8\\Multiply.scala 13:24]
  output       sign, // @[\\src\\main\\scala\\fpu8\\Multiply.scala 14:16]
  output [5:0] exponent, // @[\\src\\main\\scala\\fpu8\\Multiply.scala 15:20]
  output [2:0] fraction, // @[\\src\\main\\scala\\fpu8\\Multiply.scala 16:20]
  output       NaNFractionValue, // @[\\src\\main\\scala\\fpu8\\Multiply.scala 17:28]
  output [4:0] status // @[\\src\\main\\scala\\fpu8\\Multiply.scala 18:18]
);
  wire  _isResultNaN_T_1 = a_data[6:2] == 5'h1f; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 35:41]
  wire  _isResultNaN_T_3 = a_data[1:0] == 2'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 37:44]
  wire  _isResultNaN_T_4 = _isResultNaN_T_1 & _isResultNaN_T_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 47:24]
  wire  _isResultNaN_T_6 = b_data[6:2] == 5'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 33:39]
  wire  _isResultNaN_T_8 = b_data[1:0] == 2'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 37:44]
  wire  _isResultNaN_T_9 = _isResultNaN_T_6 & _isResultNaN_T_8; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 51:26]
  wire  _isResultNaN_T_15 = ~_isResultNaN_T_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 42:15]
  wire  _isResultNaN_T_16 = _isResultNaN_T_1 & _isResultNaN_T_15; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 41:30]
  wire  _isResultNaN_T_19 = b_data[6:2] == 5'h1f; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 35:41]
  wire  _isResultNaN_T_22 = _isResultNaN_T_19 & _isResultNaN_T_8; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 47:24]
  wire  _isResultNaN_T_24 = a_data[6:2] == 5'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 33:39]
  wire  _isResultNaN_T_27 = _isResultNaN_T_24 & _isResultNaN_T_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 51:26]
  wire  _isResultNaN_T_34 = ~_isResultNaN_T_8; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 42:15]
  wire  _isResultNaN_T_35 = _isResultNaN_T_19 & _isResultNaN_T_34; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 41:30]
  wire  isResultNaN = _isResultNaN_T_4 & _isResultNaN_T_9 | _isResultNaN_T_16 | _isResultNaN_T_22 & _isResultNaN_T_27 |
    _isResultNaN_T_35; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 443:104]
  wire  _isResultInfty_T_18 = ~_isResultNaN_T_35; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 448:62]
  wire  _isResultInfty_T_38 = ~_isResultNaN_T_16; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 448:110]
  wire  isResultInfty = _isResultNaN_T_4 & ~_isResultNaN_T_9 & ~_isResultNaN_T_35 | _isResultNaN_T_22 & ~
    _isResultNaN_T_27 & ~_isResultNaN_T_16; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 448:76]
  wire  isResult0 = _isResultNaN_T_27 & _isResultInfty_T_18 & ~_isResultNaN_T_22 | _isResultNaN_T_9 &
    _isResultInfty_T_38 & ~_isResultNaN_T_4; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 452:80]
  wire  resultNaNFractionValue = a_data[1:0] > b_data[1:0] ? a_data[0] : b_data[0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 123:18]
  wire  resultSign = a_data[7] ^ b_data[7]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 156:26]
  wire [6:0] _exponent_T_11 = {2'h0,a_data[6:2]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 168:16]
  wire [6:0] _exponent_T_13 = {2'h0,b_data[6:2]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 168:47]
  wire [6:0] _exponent_T_15 = _exponent_T_11 + _exponent_T_13; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 168:42]
  wire [6:0] _exponent_T_17 = _exponent_T_15 - 7'he; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 168:74]
  wire [6:0] _exponent_T_25 = _exponent_T_15 - 7'hf; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 169:74]
  wire [6:0] _exponent_T_26 = _isResultNaN_T_24 ^ _isResultNaN_T_6 ? _exponent_T_17 : _exponent_T_25; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 167:14]
  wire [6:0] exponent_1 = _isResultNaN_T_24 & _isResultNaN_T_6 ? 7'h1c : _exponent_T_26; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 165:12]
  wire  _firstOperandFraction_T_2 = ~_isResultNaN_T_24; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 171:36]
  wire [2:0] firstOperandFraction = {_firstOperandFraction_T_2,a_data[1:0]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 171:35]
  wire  _secondOperandFraction_T_2 = ~_isResultNaN_T_6; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 172:37]
  wire [2:0] secondOperandFraction = {_secondOperandFraction_T_2,b_data[1:0]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 172:36]
  wire [2:0] product_partialProducts_compare = secondOperandFraction[0] ? 3'h7 : 3'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 101:24]
  wire [2:0] product_partialProducts_0 = firstOperandFraction & product_partialProducts_compare; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:11]
  wire [2:0] product_partialProducts_compare_1 = secondOperandFraction[1] ? 3'h7 : 3'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 101:24]
  wire [2:0] _product_partialProducts_T_1 = firstOperandFraction & product_partialProducts_compare_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:11]
  wire [3:0] product_partialProducts_1 = {_product_partialProducts_T_1, 1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:22]
  wire [2:0] product_partialProducts_compare_2 = secondOperandFraction[2] ? 3'h7 : 3'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 101:24]
  wire [2:0] _product_partialProducts_T_2 = firstOperandFraction & product_partialProducts_compare_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:11]
  wire [4:0] product_partialProducts_2 = {_product_partialProducts_T_2, 2'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:22]
  wire [3:0] _GEN_12 = {{1'd0}, product_partialProducts_0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 112:34]
  wire [4:0] _product_partialSums_T = _GEN_12 + product_partialProducts_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 112:34]
  wire [5:0] product = _product_partialSums_T + product_partialProducts_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 112:39]
  wire [4:0] _leadingZeros_T_11 = {product[0],product[1],product[2],product[3],product[4]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 58:44]
  wire [2:0] _leadingZeros_T_17 = _leadingZeros_T_11[3] ? 3'h3 : 3'h4; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] _leadingZeros_T_18 = _leadingZeros_T_11[2] ? 3'h2 : _leadingZeros_T_17; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] _leadingZeros_T_19 = _leadingZeros_T_11[1] ? 3'h1 : _leadingZeros_T_18; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] shift = _leadingZeros_T_11[0] ? 3'h0 : _leadingZeros_T_19; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [5:0] _shiftedValue_T_3 = {product[4:0], 1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 63:23]
  wire [6:0] _shiftedValue_T_5 = {product[4:0], 2'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 63:23]
  wire [7:0] _shiftedValue_T_7 = {product[4:0], 3'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 63:23]
  wire [8:0] _shiftedValue_T_9 = {product[4:0], 4'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 63:23]
  wire [4:0] _shiftedValue_T_14 = 3'h1 == shift ? _shiftedValue_T_3[4:0] : product[4:0]; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [4:0] _shiftedValue_T_16 = 3'h2 == shift ? _shiftedValue_T_5[4:0] : _shiftedValue_T_14; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [4:0] _shiftedValue_T_18 = 3'h3 == shift ? _shiftedValue_T_7[4:0] : _shiftedValue_T_16; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [4:0] shiftedCalcValue = 3'h4 == shift ? _shiftedValue_T_9[4:0] : _shiftedValue_T_18; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [6:0] exponentShiftRight = 7'h0 - exponent_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 305:55]
  wire [6:0] exponentShiftLeft = exponent_1 - 7'h1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 308:35]
  wire  _T_2 = ~exponent_1[6]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 314:10]
  wire  _T_5 = ~exponent_1[6] & exponent_1[5:0] >= 6'h1f; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 314:40]
  wire  _T_12 = _T_2 & exponent_1[5:0] < 6'h1f; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 318:46]
  wire [4:0] _tempExponent_T_2 = exponent_1[4:0] + 5'h1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 320:38]
  wire [4:0] _tempFraction_T_3 = {product[5:2],|product[1:0]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 321:26]
  wire [5:0] _GEN_13 = {{3'd0}, shift}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 322:78]
  wire  _T_19 = _T_2 & exponent_1[5:0] > _GEN_13; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 322:46]
  wire [5:0] _tempExponent_T_5 = exponent_1[5:0] - _GEN_13; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 324:51]
  wire [4:0] _tempFraction_T_21 = 7'h0 == exponentShiftLeft ? product[4:0] : product[4:0]; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [4:0] _tempFraction_T_23 = 7'h1 == exponentShiftLeft ? _shiftedValue_T_3[4:0] : _tempFraction_T_21; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [4:0] _tempFraction_T_25 = 7'h2 == exponentShiftLeft ? _shiftedValue_T_5[4:0] : _tempFraction_T_23; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [4:0] _tempFraction_T_27 = 7'h3 == exponentShiftLeft ? _shiftedValue_T_7[4:0] : _tempFraction_T_25; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [4:0] _tempFraction_T_29 = 7'h4 == exponentShiftLeft ? _shiftedValue_T_9[4:0] : _tempFraction_T_27; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [4:0] _tempFraction_T_34 = _tempFraction_T_3 >> exponentShiftRight; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 336:110]
  wire [4:0] _GEN_0 = _T_2 & exponent_1[5:0] > 6'h0 ? _tempFraction_T_29 : _tempFraction_T_34; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 328:82 330:22 336:22]
  wire [5:0] _GEN_1 = _T_19 & shiftedCalcValue[4] ? _tempExponent_T_5 : 6'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 323:55 324:20 327:20]
  wire [4:0] _GEN_2 = _T_19 & shiftedCalcValue[4] ? shiftedCalcValue : _GEN_0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 323:55 325:20]
  wire [5:0] _GEN_3 = _T_12 & product[5] ? {{1'd0}, _tempExponent_T_2} : _GEN_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 319:54 320:20]
  wire [4:0] _GEN_4 = _T_12 & product[5] ? _tempFraction_T_3 : _GEN_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 319:54 321:20]
  wire [5:0] _GEN_5 = _T_5 & product[5] ? 6'h1f : _GEN_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 315:54 316:20]
  wire [4:0] tempFraction = _T_5 & product[5] ? 5'h1f : _GEN_4; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 315:54 317:20]
  wire  _addOne_T_2 = roundingMode == 2'h0 & tempFraction[2]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 234:42]
  wire  _addOne_T_17 = _addOne_T_2 & ~tempFraction[1] & ~tempFraction[0] & tempFraction[3]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 235:90]
  wire  _addOne_T_18 = roundingMode == 2'h0 & tempFraction[2] & (tempFraction[1] | tempFraction[0]) | _addOne_T_17; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 234:102]
  wire  _addOne_T_24 = tempFraction[2] | tempFraction[1] | tempFraction[0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 236:70]
  wire  _addOne_T_27 = roundingMode == 2'h1 & (tempFraction[2] | tempFraction[1] | tempFraction[0]) & resultSign; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 236:90]
  wire  _addOne_T_28 = _addOne_T_18 | _addOne_T_27; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 235:110]
  wire  _addOne_T_38 = roundingMode == 2'h2 & _addOne_T_24 & ~resultSign; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 237:90]
  wire  addOne = _addOne_T_28 | _addOne_T_38; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 236:106]
  wire [2:0] _GEN_15 = {{2'd0}, addOne}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 239:66]
  wire [3:0] roundedFraction = tempFraction[4:2] + _GEN_15; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 239:66]
  wire [2:0] resultFraction = roundedFraction[3] ? roundedFraction[3:1] : roundedFraction[2:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 241:28]
  wire [4:0] tempExponent = _GEN_5[4:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 310:28]
  wire [4:0] _finalExponent_T_7 = tempExponent + 5'h1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 245:20]
  wire [4:0] resultExponent = roundedFraction[3] | roundedFraction[2] & tempExponent == 5'h0 ? _finalExponent_T_7 :
    tempExponent; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 244:28]
  wire  overflow = tempExponent == 5'h1f; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 248:76]
  wire [4:0] resultStatus = {overflow,resultExponent == 5'h0,isResultNaN,isResultInfty,isResult0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 462:23]
  wire [4:0] _GEN_8 = enable ? resultExponent : 5'h0; // @[\\src\\main\\scala\\fpu8\\Multiply.scala 23:24 25:14 31:14]
  assign sign = enable & resultSign; // @[\\src\\main\\scala\\fpu8\\Multiply.scala 23:24 24:10 30:10]
  assign exponent = {{1'd0}, _GEN_8};
  assign fraction = enable ? resultFraction : 3'h0; // @[\\src\\main\\scala\\fpu8\\Multiply.scala 23:24 26:14 32:14]
  assign NaNFractionValue = enable & resultNaNFractionValue; // @[\\src\\main\\scala\\fpu8\\Multiply.scala 23:24 28:22 34:22]
  assign status = enable ? resultStatus : 5'h0; // @[\\src\\main\\scala\\fpu8\\Multiply.scala 23:24 27:12 33:12]
endmodule
module Divide(
  input        enable, // @[\\src\\main\\scala\\fpu8\\Divide.scala 10:18]
  input  [7:0] a_data, // @[\\src\\main\\scala\\fpu8\\Divide.scala 11:13]
  input  [7:0] b_data, // @[\\src\\main\\scala\\fpu8\\Divide.scala 12:13]
  input  [1:0] roundingMode, // @[\\src\\main\\scala\\fpu8\\Divide.scala 13:24]
  output       sign, // @[\\src\\main\\scala\\fpu8\\Divide.scala 14:16]
  output [5:0] exponent, // @[\\src\\main\\scala\\fpu8\\Divide.scala 15:20]
  output [2:0] fraction, // @[\\src\\main\\scala\\fpu8\\Divide.scala 16:20]
  output       NaNFractionValue, // @[\\src\\main\\scala\\fpu8\\Divide.scala 17:28]
  output [4:0] status // @[\\src\\main\\scala\\fpu8\\Divide.scala 18:18]
);
  wire  _isResultNaN_T_1 = a_data[6:2] == 5'h1f; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 35:41]
  wire  _isResultNaN_T_3 = a_data[1:0] == 2'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 37:44]
  wire  _isResultNaN_T_4 = ~_isResultNaN_T_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 42:15]
  wire  _isResultNaN_T_5 = _isResultNaN_T_1 & _isResultNaN_T_4; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 41:30]
  wire  _isResultNaN_T_7 = b_data[6:2] == 5'h1f; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 35:41]
  wire  _isResultNaN_T_9 = b_data[1:0] == 2'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 37:44]
  wire  _isResultNaN_T_10 = ~_isResultNaN_T_9; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 42:15]
  wire  _isResultNaN_T_11 = _isResultNaN_T_7 & _isResultNaN_T_10; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 41:30]
  wire  _isResultNaN_T_14 = a_data[6:2] == 5'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 33:39]
  wire  _isResultNaN_T_17 = _isResultNaN_T_14 & _isResultNaN_T_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 51:26]
  wire  _isResultNaN_T_19 = b_data[6:2] == 5'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 33:39]
  wire  _isResultNaN_T_22 = _isResultNaN_T_19 & _isResultNaN_T_9; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 51:26]
  wire  _isResultNaN_T_29 = _isResultNaN_T_1 & _isResultNaN_T_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 47:24]
  wire  _isResultNaN_T_34 = _isResultNaN_T_7 & _isResultNaN_T_9; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 47:24]
  wire  isResultNaN = _isResultNaN_T_5 | _isResultNaN_T_11 | _isResultNaN_T_17 & _isResultNaN_T_22 | _isResultNaN_T_29
     & (_isResultNaN_T_34 | _isResultNaN_T_22); // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 473:84]
  wire  _isResultInfty_T_17 = ~_isResultNaN_T_29; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 478:58]
  wire  _isResultInfty_T_25 = ~_isResultNaN_T_5; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 478:75]
  wire  _isResultInfty_T_38 = ~_isResultNaN_T_11; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 479:28]
  wire  _isResultInfty_T_45 = ~_isResultNaN_T_22; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 479:44]
  wire  _isResultInfty_T_53 = _isResultNaN_T_29 & ~_isResultNaN_T_11 & ~_isResultNaN_T_22 & ~_isResultNaN_T_34; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 479:55]
  wire  isResultInfty = _isResultNaN_T_22 & ~_isResultNaN_T_17 & ~_isResultNaN_T_29 & ~_isResultNaN_T_5 |
    _isResultInfty_T_53; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 478:88]
  wire  isResult0 = _isResultNaN_T_17 & _isResultInfty_T_45 & _isResultInfty_T_38 | _isResultNaN_T_34 &
    _isResultInfty_T_17 & _isResultInfty_T_25; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 484:72]
  wire  resultNaNFractionValue = a_data[1:0] > b_data[1:0] ? a_data[0] : b_data[0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 123:18]
  wire  resultSign = a_data[7] ^ b_data[7]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 178:26]
  wire [2:0] _tempDividendFraction_T_3 = {a_data[1:0],1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 180:10]
  wire [2:0] _tempDividendFraction_T_5 = {1'h1,a_data[1:0]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 181:10]
  wire [2:0] tempDividendFraction = _isResultNaN_T_14 ? _tempDividendFraction_T_3 : _tempDividendFraction_T_5; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 179:35]
  wire [2:0] _tempDivisorFraction_T_3 = {b_data[1:0],1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 184:10]
  wire [2:0] _tempDivisorFraction_T_5 = {1'h1,b_data[1:0]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 185:10]
  wire [2:0] tempDivisorFraction = _isResultNaN_T_19 ? _tempDivisorFraction_T_3 : _tempDivisorFraction_T_5; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 183:34]
  wire [6:0] _tempExponent_T_1 = {2'h0,a_data[6:2]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 187:27]
  wire [6:0] _tempExponent_T_3 = {2'h0,b_data[6:2]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 188:10]
  wire [6:0] _tempExponent_T_5 = _tempExponent_T_1 - _tempExponent_T_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 187:53]
  wire [6:0] tempExponent = _tempExponent_T_5 + 7'hf; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 188:37]
  wire [2:0] _leadingZeros_T_5 = {tempDividendFraction[0],tempDividendFraction[1],tempDividendFraction[2]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 58:44]
  wire [1:0] _leadingZeros_T_9 = _leadingZeros_T_5[1] ? 2'h1 : 2'h2; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [1:0] dividendShift = _leadingZeros_T_5[0] ? 2'h0 : _leadingZeros_T_9; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _shiftedValue_T_3 = {tempDividendFraction, 1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 63:23]
  wire [4:0] _shiftedValue_T_5 = {tempDividendFraction, 2'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 63:23]
  wire [2:0] _shiftedValue_T_10 = 2'h1 == dividendShift ? _shiftedValue_T_3[2:0] : tempDividendFraction; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [2:0] dividendFraction = 2'h2 == dividendShift ? _shiftedValue_T_5[2:0] : _shiftedValue_T_10; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [2:0] _leadingZeros_T_16 = {tempDivisorFraction[0],tempDivisorFraction[1],tempDivisorFraction[2]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 58:44]
  wire [1:0] _leadingZeros_T_20 = _leadingZeros_T_16[1] ? 2'h1 : 2'h2; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [1:0] divisorShift = _leadingZeros_T_16[0] ? 2'h0 : _leadingZeros_T_20; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [3:0] _shiftedValue_T_16 = {tempDivisorFraction, 1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 63:23]
  wire [4:0] _shiftedValue_T_18 = {tempDivisorFraction, 2'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 63:23]
  wire [2:0] _shiftedValue_T_23 = 2'h1 == divisorShift ? _shiftedValue_T_16[2:0] : tempDivisorFraction; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [2:0] divisorFraction = 2'h2 == divisorShift ? _shiftedValue_T_18[2:0] : _shiftedValue_T_23; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [6:0] _GEN_16 = {{5'd0}, dividendShift}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 195:33]
  wire [6:0] _exponent_T_1 = tempExponent - _GEN_16; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 195:33]
  wire [6:0] _GEN_17 = {{5'd0}, divisorShift}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 195:49]
  wire [6:0] exponent_1 = _exponent_T_1 + _GEN_17; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 195:49]
  wire [2:0] _GEN_1 = 2'h1 == divisorFraction[1:0] ? 3'h5 : 3'h7; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 203:{24,24}]
  wire [2:0] _GEN_2 = 2'h2 == divisorFraction[1:0] ? 3'h3 : _GEN_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 203:{24,24}]
  wire [2:0] _GEN_3 = 2'h3 == divisorFraction[1:0] ? 3'h1 : _GEN_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 203:{24,24}]
  wire [4:0] quotient_initGuess = {2'h1,_GEN_3}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 203:24]
  wire [4:0] quotient_secondGuess_firstStep_partialProducts_compare = divisorFraction[0] ? 5'h1f : 5'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 101:24]
  wire [4:0] quotient_secondGuess_firstStep_partialProducts_0 = quotient_initGuess &
    quotient_secondGuess_firstStep_partialProducts_compare; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:11]
  wire [4:0] quotient_secondGuess_firstStep_partialProducts_compare_1 = divisorFraction[1] ? 5'h1f : 5'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 101:24]
  wire [4:0] _quotient_secondGuess_firstStep_partialProducts_T_1 = quotient_initGuess &
    quotient_secondGuess_firstStep_partialProducts_compare_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:11]
  wire [5:0] quotient_secondGuess_firstStep_partialProducts_1 = {_quotient_secondGuess_firstStep_partialProducts_T_1
    , 1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:22]
  wire [4:0] quotient_secondGuess_firstStep_partialProducts_compare_2 = divisorFraction[2] ? 5'h1f : 5'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 101:24]
  wire [4:0] _quotient_secondGuess_firstStep_partialProducts_T_2 = quotient_initGuess &
    quotient_secondGuess_firstStep_partialProducts_compare_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:11]
  wire [6:0] quotient_secondGuess_firstStep_partialProducts_2 = {_quotient_secondGuess_firstStep_partialProducts_T_2
    , 2'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:22]
  wire [5:0] _GEN_18 = {{1'd0}, quotient_secondGuess_firstStep_partialProducts_0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 112:34]
  wire [6:0] _quotient_secondGuess_firstStep_partialSums_T = _GEN_18 + quotient_secondGuess_firstStep_partialProducts_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 112:34]
  wire [7:0] quotient_secondGuess_firstStep = _quotient_secondGuess_firstStep_partialSums_T +
    quotient_secondGuess_firstStep_partialProducts_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 112:39]
  wire [5:0] quotient_secondGuess_firstStepRnd = {1'h0,quotient_secondGuess_firstStep[6:2]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 79:12]
  wire [4:0] _quotient_secondGuess_secondStep_T_1 = ~quotient_secondGuess_firstStepRnd[4:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 214:25]
  wire [4:0] quotient_secondGuess_secondStep = _quotient_secondGuess_secondStep_T_1 + 5'h1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 214:70]
  wire [4:0] quotient_secondGuess_finalStep_partialProducts_compare = quotient_secondGuess_secondStep[0] ? 5'h1f : 5'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 101:24]
  wire [4:0] quotient_secondGuess_finalStep_partialProducts_0 = quotient_initGuess &
    quotient_secondGuess_finalStep_partialProducts_compare; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:11]
  wire [4:0] quotient_secondGuess_finalStep_partialProducts_compare_1 = quotient_secondGuess_secondStep[1] ? 5'h1f : 5'h0
    ; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 101:24]
  wire [4:0] _quotient_secondGuess_finalStep_partialProducts_T_1 = quotient_initGuess &
    quotient_secondGuess_finalStep_partialProducts_compare_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:11]
  wire [5:0] quotient_secondGuess_finalStep_partialProducts_1 = {_quotient_secondGuess_finalStep_partialProducts_T_1
    , 1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:22]
  wire [4:0] quotient_secondGuess_finalStep_partialProducts_compare_2 = quotient_secondGuess_secondStep[2] ? 5'h1f : 5'h0
    ; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 101:24]
  wire [4:0] _quotient_secondGuess_finalStep_partialProducts_T_2 = quotient_initGuess &
    quotient_secondGuess_finalStep_partialProducts_compare_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:11]
  wire [6:0] quotient_secondGuess_finalStep_partialProducts_2 = {_quotient_secondGuess_finalStep_partialProducts_T_2
    , 2'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:22]
  wire [4:0] quotient_secondGuess_finalStep_partialProducts_compare_3 = quotient_secondGuess_secondStep[3] ? 5'h1f : 5'h0
    ; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 101:24]
  wire [4:0] _quotient_secondGuess_finalStep_partialProducts_T_3 = quotient_initGuess &
    quotient_secondGuess_finalStep_partialProducts_compare_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:11]
  wire [7:0] quotient_secondGuess_finalStep_partialProducts_3 = {_quotient_secondGuess_finalStep_partialProducts_T_3
    , 3'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:22]
  wire [4:0] quotient_secondGuess_finalStep_partialProducts_compare_4 = quotient_secondGuess_secondStep[4] ? 5'h1f : 5'h0
    ; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 101:24]
  wire [4:0] _quotient_secondGuess_finalStep_partialProducts_T_4 = quotient_initGuess &
    quotient_secondGuess_finalStep_partialProducts_compare_4; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:11]
  wire [8:0] quotient_secondGuess_finalStep_partialProducts_4 = {_quotient_secondGuess_finalStep_partialProducts_T_4
    , 4'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:22]
  wire [5:0] _GEN_19 = {{1'd0}, quotient_secondGuess_finalStep_partialProducts_0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 112:34]
  wire [6:0] _quotient_secondGuess_finalStep_partialSums_T = _GEN_19 + quotient_secondGuess_finalStep_partialProducts_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 112:34]
  wire [7:0] quotient_secondGuess_finalStep_partialSums_0 = _quotient_secondGuess_finalStep_partialSums_T +
    quotient_secondGuess_finalStep_partialProducts_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 112:39]
  wire [8:0] _GEN_20 = {{1'd0}, quotient_secondGuess_finalStep_partialProducts_3}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 113:31]
  wire [9:0] quotient_secondGuess_finalStep_partialSums_1 = _GEN_20 + quotient_secondGuess_finalStep_partialProducts_4; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 113:31]
  wire [9:0] _GEN_21 = {{2'd0}, quotient_secondGuess_finalStep_partialSums_0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 109:15]
  wire [10:0] _quotient_secondGuess_finalStep_T = _GEN_21 + quotient_secondGuess_finalStep_partialSums_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 109:15]
  wire [9:0] quotient_secondGuess_finalStep = _quotient_secondGuess_finalStep_T[9:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 218:27 219:17]
  wire  _quotient_secondGuess_res_roundedValue_T_4 = quotient_secondGuess_finalStep[3] & |quotient_secondGuess_finalStep
    [2:1]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 77:59]
  wire [4:0] _GEN_22 = {{4'd0}, _quotient_secondGuess_res_roundedValue_T_4}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 77:35]
  wire [5:0] quotient_secondGuess = quotient_secondGuess_finalStep[8:4] + _GEN_22; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 77:35]
  wire [4:0] quotient_finalGuess_firstStep_partialProducts_0 = quotient_secondGuess[4:0] &
    quotient_secondGuess_firstStep_partialProducts_compare; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:11]
  wire [4:0] _quotient_finalGuess_firstStep_partialProducts_T_1 = quotient_secondGuess[4:0] &
    quotient_secondGuess_firstStep_partialProducts_compare_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:11]
  wire [5:0] quotient_finalGuess_firstStep_partialProducts_1 = {_quotient_finalGuess_firstStep_partialProducts_T_1
    , 1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:22]
  wire [4:0] _quotient_finalGuess_firstStep_partialProducts_T_2 = quotient_secondGuess[4:0] &
    quotient_secondGuess_firstStep_partialProducts_compare_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:11]
  wire [6:0] quotient_finalGuess_firstStep_partialProducts_2 = {_quotient_finalGuess_firstStep_partialProducts_T_2
    , 2'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:22]
  wire [5:0] _GEN_23 = {{1'd0}, quotient_finalGuess_firstStep_partialProducts_0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 112:34]
  wire [6:0] _quotient_finalGuess_firstStep_partialSums_T = _GEN_23 + quotient_finalGuess_firstStep_partialProducts_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 112:34]
  wire [7:0] quotient_finalGuess_firstStep = _quotient_finalGuess_firstStep_partialSums_T +
    quotient_finalGuess_firstStep_partialProducts_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 112:39]
  wire [5:0] quotient_finalGuess_firstStepRnd = {1'h0,quotient_finalGuess_firstStep[6:2]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 79:12]
  wire [4:0] _quotient_finalGuess_secondStep_T_1 = ~quotient_finalGuess_firstStepRnd[4:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 214:25]
  wire [4:0] quotient_finalGuess_secondStep = _quotient_finalGuess_secondStep_T_1 + 5'h1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 214:70]
  wire [4:0] quotient_finalGuess_finalStep_partialProducts_compare = quotient_finalGuess_secondStep[0] ? 5'h1f : 5'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 101:24]
  wire [4:0] quotient_finalGuess_finalStep_partialProducts_0 = quotient_secondGuess[4:0] &
    quotient_finalGuess_finalStep_partialProducts_compare; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:11]
  wire [4:0] quotient_finalGuess_finalStep_partialProducts_compare_1 = quotient_finalGuess_secondStep[1] ? 5'h1f : 5'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 101:24]
  wire [4:0] _quotient_finalGuess_finalStep_partialProducts_T_1 = quotient_secondGuess[4:0] &
    quotient_finalGuess_finalStep_partialProducts_compare_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:11]
  wire [5:0] quotient_finalGuess_finalStep_partialProducts_1 = {_quotient_finalGuess_finalStep_partialProducts_T_1
    , 1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:22]
  wire [4:0] quotient_finalGuess_finalStep_partialProducts_compare_2 = quotient_finalGuess_secondStep[2] ? 5'h1f : 5'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 101:24]
  wire [4:0] _quotient_finalGuess_finalStep_partialProducts_T_2 = quotient_secondGuess[4:0] &
    quotient_finalGuess_finalStep_partialProducts_compare_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:11]
  wire [6:0] quotient_finalGuess_finalStep_partialProducts_2 = {_quotient_finalGuess_finalStep_partialProducts_T_2
    , 2'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:22]
  wire [4:0] quotient_finalGuess_finalStep_partialProducts_compare_3 = quotient_finalGuess_secondStep[3] ? 5'h1f : 5'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 101:24]
  wire [4:0] _quotient_finalGuess_finalStep_partialProducts_T_3 = quotient_secondGuess[4:0] &
    quotient_finalGuess_finalStep_partialProducts_compare_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:11]
  wire [7:0] quotient_finalGuess_finalStep_partialProducts_3 = {_quotient_finalGuess_finalStep_partialProducts_T_3
    , 3'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:22]
  wire [4:0] quotient_finalGuess_finalStep_partialProducts_compare_4 = quotient_finalGuess_secondStep[4] ? 5'h1f : 5'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 101:24]
  wire [4:0] _quotient_finalGuess_finalStep_partialProducts_T_4 = quotient_secondGuess[4:0] &
    quotient_finalGuess_finalStep_partialProducts_compare_4; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:11]
  wire [8:0] quotient_finalGuess_finalStep_partialProducts_4 = {_quotient_finalGuess_finalStep_partialProducts_T_4
    , 4'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:22]
  wire [5:0] _GEN_24 = {{1'd0}, quotient_finalGuess_finalStep_partialProducts_0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 112:34]
  wire [6:0] _quotient_finalGuess_finalStep_partialSums_T = _GEN_24 + quotient_finalGuess_finalStep_partialProducts_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 112:34]
  wire [7:0] quotient_finalGuess_finalStep_partialSums_0 = _quotient_finalGuess_finalStep_partialSums_T +
    quotient_finalGuess_finalStep_partialProducts_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 112:39]
  wire [8:0] _GEN_25 = {{1'd0}, quotient_finalGuess_finalStep_partialProducts_3}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 113:31]
  wire [9:0] quotient_finalGuess_finalStep_partialSums_1 = _GEN_25 + quotient_finalGuess_finalStep_partialProducts_4; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 113:31]
  wire [9:0] _GEN_26 = {{2'd0}, quotient_finalGuess_finalStep_partialSums_0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 109:15]
  wire [10:0] _quotient_finalGuess_finalStep_T = _GEN_26 + quotient_finalGuess_finalStep_partialSums_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 109:15]
  wire [9:0] quotient_finalGuess_finalStep = _quotient_finalGuess_finalStep_T[9:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 218:27 219:17]
  wire  _quotient_finalGuess_res_roundedValue_T_4 = quotient_finalGuess_finalStep[3] & |quotient_finalGuess_finalStep[2:
    1]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 77:59]
  wire [4:0] _GEN_27 = {{4'd0}, _quotient_finalGuess_res_roundedValue_T_4}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 77:35]
  wire [5:0] quotient_finalGuess = quotient_finalGuess_finalStep[8:4] + _GEN_27; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 77:35]
  wire [4:0] quotient_partialProducts_compare = dividendFraction[0] ? 5'h1f : 5'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 101:24]
  wire [4:0] quotient_partialProducts_0 = quotient_finalGuess[4:0] & quotient_partialProducts_compare; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:11]
  wire [4:0] quotient_partialProducts_compare_1 = dividendFraction[1] ? 5'h1f : 5'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 101:24]
  wire [4:0] _quotient_partialProducts_T_1 = quotient_finalGuess[4:0] & quotient_partialProducts_compare_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:11]
  wire [5:0] quotient_partialProducts_1 = {_quotient_partialProducts_T_1, 1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:22]
  wire [4:0] quotient_partialProducts_compare_2 = dividendFraction[2] ? 5'h1f : 5'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 101:24]
  wire [4:0] _quotient_partialProducts_T_2 = quotient_finalGuess[4:0] & quotient_partialProducts_compare_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:11]
  wire [6:0] quotient_partialProducts_2 = {_quotient_partialProducts_T_2, 2'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 102:22]
  wire [5:0] _GEN_28 = {{1'd0}, quotient_partialProducts_0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 112:34]
  wire [6:0] _quotient_partialSums_T = _GEN_28 + quotient_partialProducts_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 112:34]
  wire [7:0] quotient = _quotient_partialSums_T + quotient_partialProducts_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 112:39]
  wire [6:0] _leadingZeros_T_39 = {quotient[0],quotient[1],quotient[2],quotient[3],quotient[4],quotient[5],quotient[6]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 58:44]
  wire [2:0] _leadingZeros_T_47 = _leadingZeros_T_39[5] ? 3'h5 : 3'h6; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] _leadingZeros_T_48 = _leadingZeros_T_39[4] ? 3'h4 : _leadingZeros_T_47; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] _leadingZeros_T_49 = _leadingZeros_T_39[3] ? 3'h3 : _leadingZeros_T_48; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] _leadingZeros_T_50 = _leadingZeros_T_39[2] ? 3'h2 : _leadingZeros_T_49; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] _leadingZeros_T_51 = _leadingZeros_T_39[1] ? 3'h1 : _leadingZeros_T_50; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [2:0] shift = _leadingZeros_T_39[0] ? 3'h0 : _leadingZeros_T_51; // @[src/main/scala/chisel3/util/Mux.scala 50:70]
  wire [7:0] _shiftedValue_T_29 = {quotient[6:0], 1'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 63:23]
  wire [8:0] _shiftedValue_T_31 = {quotient[6:0], 2'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 63:23]
  wire [9:0] _shiftedValue_T_33 = {quotient[6:0], 3'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 63:23]
  wire [10:0] _shiftedValue_T_35 = {quotient[6:0], 4'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 63:23]
  wire [11:0] _shiftedValue_T_37 = {quotient[6:0], 5'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 63:23]
  wire [12:0] _shiftedValue_T_39 = {quotient[6:0], 6'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 63:23]
  wire [6:0] _shiftedValue_T_44 = 3'h1 == shift ? _shiftedValue_T_29[6:0] : quotient[6:0]; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [6:0] _shiftedValue_T_46 = 3'h2 == shift ? _shiftedValue_T_31[6:0] : _shiftedValue_T_44; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [6:0] _shiftedValue_T_48 = 3'h3 == shift ? _shiftedValue_T_33[6:0] : _shiftedValue_T_46; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [6:0] _shiftedValue_T_50 = 3'h4 == shift ? _shiftedValue_T_35[6:0] : _shiftedValue_T_48; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [6:0] _shiftedValue_T_52 = 3'h5 == shift ? _shiftedValue_T_37[6:0] : _shiftedValue_T_50; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [6:0] shiftedCalcValue = 3'h6 == shift ? _shiftedValue_T_39[6:0] : _shiftedValue_T_52; // @[src/main/scala/chisel3/util/Mux.scala 77:13]
  wire [6:0] exponentShiftRight = 7'h0 - exponent_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 352:55]
  wire [6:0] exponentShiftLeft = exponent_1 - 7'h1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 355:35]
  wire  _T_2 = ~exponent_1[6]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 363:10]
  wire  _T_5 = ~exponent_1[6] & exponent_1[5:0] >= 6'h1f; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 363:40]
  wire  _T_12 = _T_2 & exponent_1[5:0] < 6'h1f; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 367:46]
  wire [5:0] _tempExponent_T_9 = exponent_1[5:0] + 6'h1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 369:51]
  wire [5:0] _GEN_29 = {{3'd0}, shift}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 377:78]
  wire  _T_19 = _T_2 & exponent_1[5:0] > _GEN_29; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 377:46]
  wire [5:0] _tempExponent_T_12 = exponent_1[5:0] - _GEN_29; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 379:51]
  wire [132:0] _GEN_0 = {{127'd0}, quotient[6:1]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 395:83]
  wire [132:0] _tempFraction_T_3 = _GEN_0 << exponentShiftLeft; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 395:83]
  wire  _tempFraction_T_6 = &quotient[1:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 399:125]
  wire [5:0] _GEN_31 = {{5'd0}, _tempFraction_T_6}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 398:118]
  wire [5:0] _tempFraction_T_8 = quotient[7:2] + _GEN_31; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 398:118]
  wire [5:0] _tempFraction_T_9 = _tempFraction_T_8 >> exponentShiftRight; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 399:138]
  wire [132:0] _GEN_4 = _T_2 & exponent_1[5:0] > 6'h0 ? _tempFraction_T_3 : {{127'd0}, _tempFraction_T_9}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 389:82 390:22 398:22]
  wire [5:0] _GEN_5 = _T_19 & shiftedCalcValue[6] ? _tempExponent_T_12 : 6'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 378:55 379:20 388:20]
  wire [132:0] _GEN_6 = _T_19 & shiftedCalcValue[6] ? {{127'd0}, shiftedCalcValue[6:1]} : _GEN_4; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 378:55 380:20]
  wire [5:0] _GEN_7 = _T_12 & quotient[7] ? _tempExponent_T_9 : _GEN_5; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 368:54 369:20]
  wire [132:0] _GEN_8 = _T_12 & quotient[7] ? {{127'd0}, quotient[6:1]} : _GEN_6; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 368:54 370:20]
  wire [5:0] tempExponent_1 = _T_5 & quotient[7] ? 6'h1f : _GEN_7; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 364:54 365:20]
  wire [132:0] _GEN_10 = _T_5 & quotient[7] ? 133'h7f : _GEN_8; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 364:54 366:20]
  wire [6:0] tempFraction = _GEN_10[6:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 359:28]
  wire  _addOne_T_2 = roundingMode == 2'h0 & tempFraction[2]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 234:42]
  wire  _addOne_T_17 = _addOne_T_2 & ~tempFraction[1] & ~tempFraction[0] & tempFraction[3]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 235:90]
  wire  _addOne_T_18 = roundingMode == 2'h0 & tempFraction[2] & (tempFraction[1] | tempFraction[0]) | _addOne_T_17; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 234:102]
  wire  _addOne_T_24 = tempFraction[2] | tempFraction[1] | tempFraction[0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 236:70]
  wire  _addOne_T_27 = roundingMode == 2'h1 & (tempFraction[2] | tempFraction[1] | tempFraction[0]) & resultSign; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 236:90]
  wire  _addOne_T_28 = _addOne_T_18 | _addOne_T_27; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 235:110]
  wire  _addOne_T_38 = roundingMode == 2'h2 & _addOne_T_24 & ~resultSign; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 237:90]
  wire  addOne = _addOne_T_28 | _addOne_T_38; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 236:106]
  wire [2:0] _GEN_32 = {{2'd0}, addOne}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 239:66]
  wire [3:0] roundedFraction = tempFraction[5:3] + _GEN_32; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 239:66]
  wire [2:0] resultFraction = roundedFraction[3] ? roundedFraction[3:1] : roundedFraction[2:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 241:28]
  wire [5:0] _finalExponent_T_7 = tempExponent_1 + 6'h1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 245:20]
  wire [5:0] resultExponent = roundedFraction[3] | roundedFraction[2] & tempExponent_1 == 6'h0 ? _finalExponent_T_7 :
    tempExponent_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 244:28]
  wire  overflow = resultExponent >= 6'h20 | tempExponent_1 == 6'h1f; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 248:59]
  wire [4:0] resultStatus = {overflow,resultExponent == 6'h0,isResultNaN,isResultInfty,isResult0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 496:23]
  assign sign = enable & resultSign; // @[\\src\\main\\scala\\fpu8\\Divide.scala 23:24 24:10 30:10]
  assign exponent = enable ? resultExponent : 6'h0; // @[\\src\\main\\scala\\fpu8\\Divide.scala 23:24 25:14 31:14]
  assign fraction = enable ? resultFraction : 3'h0; // @[\\src\\main\\scala\\fpu8\\Divide.scala 23:24 26:14 32:14]
  assign NaNFractionValue = enable & resultNaNFractionValue; // @[\\src\\main\\scala\\fpu8\\Divide.scala 23:24 28:22 34:22]
  assign status = enable ? resultStatus : 5'h0; // @[\\src\\main\\scala\\fpu8\\Divide.scala 23:24 27:12 33:12]
endmodule
module Compare(
  input        enable, // @[\\src\\main\\scala\\fpu8\\Compare.scala 6:18]
  input  [2:0] compareMode, // @[\\src\\main\\scala\\fpu8\\Compare.scala 7:23]
  input  [7:0] a_data, // @[\\src\\main\\scala\\fpu8\\Compare.scala 8:13]
  input  [7:0] b_data, // @[\\src\\main\\scala\\fpu8\\Compare.scala 9:13]
  output [7:0] z, // @[\\src\\main\\scala\\fpu8\\Compare.scala 10:13]
  output [4:0] status // @[\\src\\main\\scala\\fpu8\\Compare.scala 11:18]
);
  wire  _result_T_7 = a_data[6:0] > b_data[6:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 29:77]
  wire  _result_T_11 = ~a_data[7]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 506:96]
  wire  _result_T_15 = ~_result_T_7; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 506:107]
  wire [7:0] result_result = a_data[7] > b_data[7] | a_data[7] & _result_T_7 | ~a_data[7] & ~_result_T_7 ? 8'h3c : 8'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 506:132 508:14 510:14]
  wire [7:0] result_result_1 = a_data[7] < b_data[7] | a_data[7] & _result_T_15 | _result_T_11 & _result_T_7 ? 8'h3c : 8'h0
    ; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 519:133 521:14 523:14]
  wire [7:0] result_result_2 = a_data == b_data ? 8'h3c : 8'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 532:36 534:14 536:14]
  wire [7:0] _result_T_56 = result_result ^ result_result_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 544:20]
  wire [7:0] _result_T_76 = result_result_1 ^ result_result_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 550:20]
  wire  _T_6 = compareMode == 3'h5; // @[\\src\\main\\scala\\fpu8\\Compare.scala 27:28]
  wire  _result_T_79 = a_data[6:2] == 5'h1f; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 35:41]
  wire  _result_T_81 = a_data[1:0] == 2'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 37:44]
  wire  _result_T_82 = ~_result_T_81; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 42:15]
  wire  _result_T_83 = _result_T_79 & _result_T_82; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 41:30]
  wire  _result_T_85 = b_data[6:2] == 5'h1f; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 35:41]
  wire  _result_T_87 = b_data[1:0] == 2'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 37:44]
  wire  _result_T_88 = ~_result_T_87; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 42:15]
  wire  _result_T_89 = _result_T_85 & _result_T_88; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 41:30]
  wire [7:0] result_result_7 = a_data != b_data | _result_T_83 & _result_T_89 ? 8'h3c : 8'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 557:69 559:14 561:14]
  wire [7:0] _GEN_8 = compareMode == 3'h5 ? result_result_7 : 8'h0; // @[\\src\\main\\scala\\fpu8\\Compare.scala 27:36 28:14 30:14]
  wire [7:0] _GEN_9 = compareMode == 3'h4 ? _result_T_76 : _GEN_8; // @[\\src\\main\\scala\\fpu8\\Compare.scala 25:37 26:14]
  wire [7:0] _GEN_10 = compareMode == 3'h3 ? _result_T_56 : _GEN_9; // @[\\src\\main\\scala\\fpu8\\Compare.scala 23:37 24:14]
  wire [7:0] _GEN_11 = compareMode == 3'h2 ? result_result_2 : _GEN_10; // @[\\src\\main\\scala\\fpu8\\Compare.scala 21:37 22:14]
  wire [7:0] _GEN_12 = compareMode == 3'h1 ? result_result_1 : _GEN_11; // @[\\src\\main\\scala\\fpu8\\Compare.scala 19:37 20:14]
  wire [7:0] _GEN_13 = compareMode == 3'h0 ? result_result : _GEN_12; // @[\\src\\main\\scala\\fpu8\\Compare.scala 17:31 18:14]
  wire [7:0] result = enable ? _GEN_13 : 8'h0; // @[\\src\\main\\scala\\fpu8\\Compare.scala 16:23 43:12]
  wire [7:0] _z_T_15 = _T_6 & _result_T_83 & _result_T_89 ? result : 8'h0; // @[\\src\\main\\scala\\fpu8\\Compare.scala 37:15]
  wire  isNaN = enable & (_result_T_83 | _result_T_89); // @[\\src\\main\\scala\\fpu8\\Compare.scala 16:23 33:11 45:11]
  wire [2:0] _GEN_14 = isNaN ? 3'h4 : 3'h0; // @[\\src\\main\\scala\\fpu8\\Compare.scala 35:16 36:14 39:14]
  wire [7:0] _GEN_15 = isNaN ? _z_T_15 : result; // @[\\src\\main\\scala\\fpu8\\Compare.scala 35:16 37:9 40:9]
  wire [2:0] _GEN_18 = enable ? _GEN_14 : 3'h0; // @[\\src\\main\\scala\\fpu8\\Compare.scala 16:23 46:12]
  assign z = enable ? _GEN_15 : 8'h0; // @[\\src\\main\\scala\\fpu8\\Compare.scala 16:23 44:7]
  assign status = {{2'd0}, _GEN_18};
endmodule
module Convert(
  input        enable, // @[\\src\\main\\scala\\fpu8\\Convert.scala 6:18]
  input  [7:0] a_data, // @[\\src\\main\\scala\\fpu8\\Convert.scala 7:13]
  input  [1:0] roundingMode, // @[\\src\\main\\scala\\fpu8\\Convert.scala 8:24]
  input        saturationMode, // @[\\src\\main\\scala\\fpu8\\Convert.scala 9:26]
  output [7:0] z, // @[\\src\\main\\scala\\fpu8\\Convert.scala 10:13]
  output [4:0] status // @[\\src\\main\\scala\\fpu8\\Convert.scala 11:18]
);
  wire  _isResultNaN_T_1 = a_data[6:2] == 5'h1f; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 35:41]
  wire  _isResultNaN_T_3 = a_data[1:0] == 2'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 37:44]
  wire  _isResultNaN_T_4 = ~_isResultNaN_T_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 42:15]
  wire  _isResultNaN_T_5 = _isResultNaN_T_1 & _isResultNaN_T_4; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 41:30]
  wire  _isResultNaN_T_10 = _isResultNaN_T_1 & _isResultNaN_T_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 47:24]
  wire  isResultNaN = _isResultNaN_T_5 | _isResultNaN_T_10; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 605:29]
  wire  _fraction_T_1 = a_data[6:2] == 5'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 33:39]
  wire  _fraction_T_2 = ~_fraction_T_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 607:24]
  wire [5:0] tempExponent = a_data[6:2] - 5'h8; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 609:33]
  wire  isDenormalized = tempExponent[5] | tempExponent[4:0] == 5'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 611:55]
  wire  overflow = ~tempExponent[5] & tempExponent[4]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 612:50]
  wire [6:0] _shift_T = 6'h1 - tempExponent; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 613:41]
  wire [6:0] shift = isDenormalized ? _shift_T : 7'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 613:20]
  wire [6:0] _tempFraction_T = {_fraction_T_2,a_data[1:0],4'h0}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 615:27]
  wire [6:0] tempFraction = _tempFraction_T >> shift; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 615:67]
  wire  _addOne_T = roundingMode == 2'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 617:33]
  wire  _addOne_T_2 = roundingMode == 2'h0 & tempFraction[2]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 617:42]
  wire  _addOne_T_17 = _addOne_T_2 & ~tempFraction[1] & ~tempFraction[0] & tempFraction[3]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 618:90]
  wire  _addOne_T_18 = roundingMode == 2'h0 & tempFraction[2] & (tempFraction[1] | tempFraction[0]) | _addOne_T_17; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 617:102]
  wire  _addOne_T_19 = roundingMode == 2'h1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 619:22]
  wire  _addOne_T_24 = tempFraction[2] | tempFraction[1] | tempFraction[0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 619:70]
  wire  _addOne_T_28 = roundingMode == 2'h1 & (tempFraction[2] | tempFraction[1] | tempFraction[0]) & a_data[7]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 619:90]
  wire  _addOne_T_29 = _addOne_T_18 | _addOne_T_28; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 618:110]
  wire  _addOne_T_30 = roundingMode == 2'h2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 620:22]
  wire  _addOne_T_39 = ~a_data[7]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 620:93]
  wire  _addOne_T_40 = roundingMode == 2'h2 & _addOne_T_24 & ~a_data[7]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 620:90]
  wire  addOne = _addOne_T_29 | _addOne_T_40; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 619:106]
  wire [3:0] _GEN_9 = {{3'd0}, addOne}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 622:80]
  wire [4:0] roundedFraction = tempFraction[6:3] + _GEN_9; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 622:80]
  wire [3:0] _finalExponent_T_1 = isDenormalized ? 4'h0 : tempExponent[3:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 625:10]
  wire [3:0] finalExponent = overflow ? 4'hf : _finalExponent_T_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 624:28]
  wire [3:0] finalFraction = roundedFraction[3:0]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 627:40]
  wire  _T_3 = ~saturationMode; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 634:54]
  wire  _T_10 = _addOne_T_19 & _T_3 & _addOne_T_39; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 635:59]
  wire  _T_11 = _addOne_T & ~saturationMode | _T_10; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 634:63]
  wire  _T_17 = _addOne_T_30 & _T_3 & _addOne_T_39; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 636:59]
  wire  _T_18 = _T_11 | _T_17; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 635:76]
  wire  _T_24 = roundingMode == 2'h3 & _T_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 639:33]
  wire  _T_25 = _addOne_T & saturationMode | _T_24; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 638:69]
  wire [7:0] _result_T_2 = {a_data[7],4'hf,3'h6}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 640:24]
  wire  _T_35 = _addOne_T_30 & a_data[7]; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 642:33]
  wire  _T_36 = _addOne_T_19 & saturationMode & _addOne_T_39 | _T_35; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 641:85]
  wire  _T_46 = _addOne_T_30 & saturationMode & _addOne_T_39; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 645:59]
  wire  _T_47 = _addOne_T_19 & a_data[7] | _T_46; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 644:59]
  wire [7:0] _GEN_0 = _T_47 ? _result_T_2 : 8'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 645:77 646:18 648:18]
  wire [7:0] _GEN_1 = _T_36 ? _result_T_2 : _GEN_0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 642:51 643:18]
  wire [7:0] _GEN_2 = _T_25 ? _result_T_2 : _GEN_1; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 639:61 640:18]
  wire [7:0] _GEN_3 = _T_18 ? 8'h7f : _GEN_2; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 636:77 637:18]
  wire [7:0] _result_T_9 = {a_data[7],finalExponent,finalFraction[2:0]}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 651:22]
  wire [7:0] _GEN_4 = overflow ? _GEN_3 : _result_T_9; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 633:22 651:16]
  wire [7:0] _GEN_5 = isResultNaN ? 8'h7f : 8'h0; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 653:29 654:14 656:14]
  wire [7:0] result = ~isResultNaN ? _GEN_4 : _GEN_5; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 632:24]
  wire  _status_T_4 = _fraction_T_1 & _isResultNaN_T_3; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 51:26]
  wire [4:0] resultStatus = {overflow,isDenormalized,isResultNaN,1'h0,_status_T_4}; // @[\\src\\main\\scala\\fpu8\\FloatingPoint.scala 658:18]
  assign z = enable ? result : 8'h0; // @[\\src\\main\\scala\\fpu8\\Convert.scala 13:23 19:7 22:7]
  assign status = enable ? resultStatus : 5'h0; // @[\\src\\main\\scala\\fpu8\\Convert.scala 13:23 20:12 23:12]
endmodule
module GenerateFinalResult(
  input        enable, // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 12:18]
  input        sign, // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 13:16]
  input  [4:0] exponent, // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 14:20]
  input  [1:0] mantissa, // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 15:20]
  input  [1:0] roundingMode, // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 16:24]
  input        overflow, // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 17:20]
  input        saturationMode, // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 18:26]
  input        isInfty, // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 19:19]
  input        is0, // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 20:15]
  input        isNaN, // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 21:17]
  input        NaNFractionValue, // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 22:28]
  output [7:0] z // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 23:13]
);
  wire  _result_T_4 = ~isInfty; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 70:10]
  wire  _result_T_5 = ~is0; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 70:22]
  wire  _result_T_7 = ~isNaN; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 70:30]
  wire  _result_T_9 = roundingMode == 2'h0; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 72:27]
  wire  _result_T_10 = ~saturationMode; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 72:53]
  wire [7:0] _result_z_T = {sign,5'h1f,2'h0}; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 73:19]
  wire [7:0] _result_z_T_1 = {sign,5'h1e,2'h3}; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 75:19]
  wire  _result_T_17 = roundingMode == 2'h1; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 76:33]
  wire  _result_T_20 = ~sign; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 76:75]
  wire  _result_T_27 = roundingMode == 2'h2; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 78:102]
  wire [7:0] _GEN_0 = _result_T_27 & _result_T_10 & _result_T_20 ? 8'h7c : 8'h0; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 82:84 83:13 85:13]
  wire [7:0] _GEN_1 = _result_T_17 & sign | _result_T_27 & saturationMode & _result_T_20 ? 8'h7b : _GEN_0; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 80:128 81:13]
  wire [7:0] _GEN_2 = _result_T_17 & saturationMode & _result_T_20 | roundingMode == 2'h2 & sign ? 8'hfb : _GEN_1; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 78:128 79:13]
  wire [7:0] _GEN_3 = roundingMode == 2'h1 & _result_T_10 & ~sign ? 8'hfc : _GEN_2; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 76:84 77:13]
  wire [7:0] _GEN_4 = _result_T_9 & saturationMode | roundingMode == 2'h3 ? _result_z_T_1 : _GEN_3; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 74:94 75:13]
  wire [7:0] _GEN_5 = roundingMode == 2'h0 & ~saturationMode ? _result_z_T : _GEN_4; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 72:62 73:13]
  wire [7:0] _result_z_T_6 = {sign,exponent,mantissa}; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 88:17]
  wire [7:0] _GEN_6 = overflow ? _GEN_5 : _result_z_T_6; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 71:22 88:11]
  wire [7:0] _result_z_T_8 = {sign,5'h0,2'h0}; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 93:15]
  wire [7:0] _result_z_T_9 = {6'h1f,1'h1,NaNFractionValue}; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 95:15]
  wire [7:0] _GEN_7 = isNaN ? _result_z_T_9 : 8'h0; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 94:23 95:9 97:9]
  wire [7:0] _GEN_8 = _result_T_4 & is0 & _result_T_7 ? _result_z_T_8 : _GEN_7; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 92:43 93:9]
  wire [7:0] _GEN_9 = isInfty & _result_T_5 & _result_T_7 ? _result_z_T : _GEN_8; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 90:43 91:9]
  wire [7:0] result = ~isInfty & ~is0 & ~isNaN ? _GEN_6 : _GEN_9; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 70:38]
  assign z = enable ? result : 8'h0; // @[\\src\\main\\scala\\fpu8\\GenerateFinalResult.scala 31:23 32:7 34:7]
endmodule
module FPU8Generator(
  input        clock,
  input        reset,
  input        enable, // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 9:18]
  input  [7:0] a_data, // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 10:13]
  input  [7:0] b_data, // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 11:13]
  input  [3:0] opCode, // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 12:18]
  input  [1:0] roundingMode, // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 13:24]
  input        saturationMode, // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 14:26]
  output [7:0] z, // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 15:13]
  output [4:0] status // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 16:18]
);
  wire  addSub_enable; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 18:22]
  wire [7:0] addSub_a_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 18:22]
  wire [7:0] addSub_b_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 18:22]
  wire  addSub_subtract; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 18:22]
  wire [1:0] addSub_roundingMode; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 18:22]
  wire  addSub_sign; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 18:22]
  wire [5:0] addSub_exponent; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 18:22]
  wire [2:0] addSub_fraction; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 18:22]
  wire  addSub_NaNFractionValue; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 18:22]
  wire [4:0] addSub_status; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 18:22]
  wire  multiply_enable; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 20:24]
  wire [7:0] multiply_a_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 20:24]
  wire [7:0] multiply_b_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 20:24]
  wire [1:0] multiply_roundingMode; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 20:24]
  wire  multiply_sign; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 20:24]
  wire [5:0] multiply_exponent; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 20:24]
  wire [2:0] multiply_fraction; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 20:24]
  wire  multiply_NaNFractionValue; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 20:24]
  wire [4:0] multiply_status; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 20:24]
  wire  divide_enable; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 22:22]
  wire [7:0] divide_a_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 22:22]
  wire [7:0] divide_b_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 22:22]
  wire [1:0] divide_roundingMode; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 22:22]
  wire  divide_sign; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 22:22]
  wire [5:0] divide_exponent; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 22:22]
  wire [2:0] divide_fraction; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 22:22]
  wire  divide_NaNFractionValue; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 22:22]
  wire [4:0] divide_status; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 22:22]
  wire  compare_enable; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 24:23]
  wire [2:0] compare_compareMode; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 24:23]
  wire [7:0] compare_a_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 24:23]
  wire [7:0] compare_b_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 24:23]
  wire [7:0] compare_z; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 24:23]
  wire [4:0] compare_status; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 24:23]
  wire  convert_enable; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 26:23]
  wire [7:0] convert_a_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 26:23]
  wire [1:0] convert_roundingMode; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 26:23]
  wire  convert_saturationMode; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 26:23]
  wire [7:0] convert_z; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 26:23]
  wire [4:0] convert_status; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 26:23]
  wire  generateFinalResult_enable; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 28:35]
  wire  generateFinalResult_sign; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 28:35]
  wire [4:0] generateFinalResult_exponent; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 28:35]
  wire [1:0] generateFinalResult_mantissa; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 28:35]
  wire [1:0] generateFinalResult_roundingMode; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 28:35]
  wire  generateFinalResult_overflow; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 28:35]
  wire  generateFinalResult_saturationMode; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 28:35]
  wire  generateFinalResult_isInfty; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 28:35]
  wire  generateFinalResult_is0; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 28:35]
  wire  generateFinalResult_isNaN; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 28:35]
  wire  generateFinalResult_NaNFractionValue; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 28:35]
  wire [7:0] generateFinalResult_z; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 28:35]
  wire  _addSub_enable_T_2 = opCode == 4'h0 | opCode == 4'h1; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 30:39]
  wire  _multiply_enable_T = opCode == 4'h2; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 36:33]
  wire  _divide_enable_T = opCode == 4'h3; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 41:31]
  wire  _compare_enable_T = opCode == 4'h4; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 46:32]
  wire  _compare_enable_T_1 = opCode == 4'h5; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 46:50]
  wire  _compare_enable_T_3 = opCode == 4'h6; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 46:68]
  wire  _compare_enable_T_5 = opCode == 4'h7; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 46:86]
  wire  _compare_enable_T_7 = opCode == 4'h8; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 46:104]
  wire  _compare_enable_T_10 = opCode == 4'h4 | opCode == 4'h5 | opCode == 4'h6 | opCode == 4'h7 | opCode == 4'h8 |
    opCode == 4'h9; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 46:112]
  wire [2:0] _compare_compareMode_T_5 = _compare_enable_T_7 ? 3'h4 : 3'h5; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 52:14]
  wire [2:0] _compare_compareMode_T_6 = _compare_enable_T_5 ? 3'h3 : _compare_compareMode_T_5; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 51:12]
  wire [2:0] _compare_compareMode_T_7 = _compare_enable_T_3 ? 3'h2 : _compare_compareMode_T_6; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 50:10]
  wire [2:0] _compare_compareMode_T_8 = _compare_enable_T_1 ? 3'h1 : _compare_compareMode_T_7; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 49:8]
  wire  _convert_enable_T = opCode == 4'ha; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 56:32]
  wire [7:0] _GEN_1 = _convert_enable_T ? convert_z : 8'h0; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 119:30 131:7 145:7]
  wire [4:0] _GEN_2 = _convert_enable_T ? convert_status : 5'h0; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 119:30 132:12 146:12]
  wire [7:0] _GEN_4 = _compare_enable_T_10 ? compare_z : _GEN_1; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 105:119 117:7]
  wire [4:0] _GEN_5 = _compare_enable_T_10 ? compare_status : _GEN_2; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 105:119 118:12]
  wire  _GEN_6 = _divide_enable_T & divide_sign; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 91:30 92:30]
  wire [4:0] _GEN_7 = _divide_enable_T ? divide_exponent[4:0] : 5'h0; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 91:30 93:34]
  wire [1:0] _GEN_8 = _divide_enable_T ? divide_fraction[1:0] : 2'h0; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 91:30 94:34]
  wire [1:0] _GEN_9 = _divide_enable_T ? roundingMode : 2'h0; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 91:30 95:38]
  wire  _GEN_10 = _divide_enable_T & divide_status[4]; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 91:30 96:34]
  wire  _GEN_11 = _divide_enable_T & saturationMode; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 91:30 97:40]
  wire  _GEN_12 = _divide_enable_T & divide_status[1]; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 91:30 98:33]
  wire  _GEN_13 = _divide_enable_T & divide_status[0]; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 91:30 99:29]
  wire  _GEN_14 = _divide_enable_T & divide_status[2]; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 91:30 100:31]
  wire  _GEN_15 = _divide_enable_T & divide_NaNFractionValue; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 91:30 101:42]
  wire [7:0] _GEN_16 = _divide_enable_T ? generateFinalResult_z : _GEN_4; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 91:30 103:7]
  wire [4:0] _GEN_17 = _divide_enable_T ? divide_status : _GEN_5; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 104:12 91:30]
  wire  _GEN_18 = _multiply_enable_T ? multiply_sign : _GEN_6; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 77:30 78:30]
  wire [4:0] _GEN_19 = _multiply_enable_T ? multiply_exponent[4:0] : _GEN_7; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 77:30 79:34]
  wire [1:0] _GEN_20 = _multiply_enable_T ? multiply_fraction[1:0] : _GEN_8; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 77:30 80:34]
  wire [1:0] _GEN_21 = _multiply_enable_T ? roundingMode : _GEN_9; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 77:30 81:38]
  wire  _GEN_22 = _multiply_enable_T ? multiply_status[4] : _GEN_10; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 77:30 82:34]
  wire  _GEN_23 = _multiply_enable_T ? saturationMode : _GEN_11; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 77:30 83:40]
  wire  _GEN_24 = _multiply_enable_T ? multiply_status[1] : _GEN_12; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 77:30 84:33]
  wire  _GEN_25 = _multiply_enable_T ? multiply_status[0] : _GEN_13; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 77:30 85:29]
  wire  _GEN_26 = _multiply_enable_T ? multiply_status[2] : _GEN_14; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 77:30 86:31]
  wire  _GEN_27 = _multiply_enable_T ? multiply_NaNFractionValue : _GEN_15; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 77:30 87:42]
  wire [7:0] _GEN_28 = _multiply_enable_T ? generateFinalResult_z : _GEN_16; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 77:30 89:7]
  wire [4:0] _GEN_29 = _multiply_enable_T ? multiply_status : _GEN_17; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 77:30 90:12]
  Add addSub ( // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 18:22]
    .enable(addSub_enable),
    .a_data(addSub_a_data),
    .b_data(addSub_b_data),
    .subtract(addSub_subtract),
    .roundingMode(addSub_roundingMode),
    .sign(addSub_sign),
    .exponent(addSub_exponent),
    .fraction(addSub_fraction),
    .NaNFractionValue(addSub_NaNFractionValue),
    .status(addSub_status)
  );
  Multiply multiply ( // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 20:24]
    .enable(multiply_enable),
    .a_data(multiply_a_data),
    .b_data(multiply_b_data),
    .roundingMode(multiply_roundingMode),
    .sign(multiply_sign),
    .exponent(multiply_exponent),
    .fraction(multiply_fraction),
    .NaNFractionValue(multiply_NaNFractionValue),
    .status(multiply_status)
  );
  Divide divide ( // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 22:22]
    .enable(divide_enable),
    .a_data(divide_a_data),
    .b_data(divide_b_data),
    .roundingMode(divide_roundingMode),
    .sign(divide_sign),
    .exponent(divide_exponent),
    .fraction(divide_fraction),
    .NaNFractionValue(divide_NaNFractionValue),
    .status(divide_status)
  );
  Compare compare ( // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 24:23]
    .enable(compare_enable),
    .compareMode(compare_compareMode),
    .a_data(compare_a_data),
    .b_data(compare_b_data),
    .z(compare_z),
    .status(compare_status)
  );
  Convert convert ( // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 26:23]
    .enable(convert_enable),
    .a_data(convert_a_data),
    .roundingMode(convert_roundingMode),
    .saturationMode(convert_saturationMode),
    .z(convert_z),
    .status(convert_status)
  );
  GenerateFinalResult generateFinalResult ( // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 28:35]
    .enable(generateFinalResult_enable),
    .sign(generateFinalResult_sign),
    .exponent(generateFinalResult_exponent),
    .mantissa(generateFinalResult_mantissa),
    .roundingMode(generateFinalResult_roundingMode),
    .overflow(generateFinalResult_overflow),
    .saturationMode(generateFinalResult_saturationMode),
    .isInfty(generateFinalResult_isInfty),
    .is0(generateFinalResult_is0),
    .isNaN(generateFinalResult_isNaN),
    .NaNFractionValue(generateFinalResult_NaNFractionValue),
    .z(generateFinalResult_z)
  );
  assign z = _addSub_enable_T_2 ? generateFinalResult_z : _GEN_28; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 63:42 75:7]
  assign status = _addSub_enable_T_2 ? addSub_status : _GEN_29; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 63:42 76:12]
  assign addSub_enable = (opCode == 4'h0 | opCode == 4'h1) & enable; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 30:23]
  assign addSub_a_data = a_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 31:12]
  assign addSub_b_data = b_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 32:12]
  assign addSub_subtract = opCode == 4'h1; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 33:33]
  assign addSub_roundingMode = roundingMode; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 34:23]
  assign multiply_enable = opCode == 4'h2 & enable; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 36:25]
  assign multiply_a_data = a_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 37:14]
  assign multiply_b_data = b_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 38:14]
  assign multiply_roundingMode = roundingMode; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 39:25]
  assign divide_enable = opCode == 4'h3 & enable; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 41:23]
  assign divide_a_data = a_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 42:12]
  assign divide_b_data = b_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 43:12]
  assign divide_roundingMode = roundingMode; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 44:23]
  assign compare_enable = (opCode == 4'h4 | opCode == 4'h5 | opCode == 4'h6 | opCode == 4'h7 | opCode == 4'h8 | opCode
     == 4'h9) & enable; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 46:24]
  assign compare_compareMode = _compare_enable_T ? 3'h0 : _compare_compareMode_T_8; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 48:29]
  assign compare_a_data = a_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 53:13]
  assign compare_b_data = b_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 54:13]
  assign convert_enable = opCode == 4'ha & enable; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 56:24]
  assign convert_a_data = a_data; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 57:13]
  assign convert_roundingMode = roundingMode; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 58:24]
  assign convert_saturationMode = saturationMode; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 59:26]
  assign generateFinalResult_enable = enable; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 61:30]
  assign generateFinalResult_sign = _addSub_enable_T_2 ? addSub_sign : _GEN_18; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 63:42 64:30]
  assign generateFinalResult_exponent = _addSub_enable_T_2 ? addSub_exponent[4:0] : _GEN_19; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 63:42 65:34]
  assign generateFinalResult_mantissa = _addSub_enable_T_2 ? addSub_fraction[1:0] : _GEN_20; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 63:42 66:34]
  assign generateFinalResult_roundingMode = _addSub_enable_T_2 ? roundingMode : _GEN_21; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 63:42 67:38]
  assign generateFinalResult_overflow = _addSub_enable_T_2 ? addSub_status[4] : _GEN_22; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 63:42 68:34]
  assign generateFinalResult_saturationMode = _addSub_enable_T_2 ? saturationMode : _GEN_23; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 63:42 69:40]
  assign generateFinalResult_isInfty = _addSub_enable_T_2 ? addSub_status[1] : _GEN_24; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 63:42 70:33]
  assign generateFinalResult_is0 = _addSub_enable_T_2 ? addSub_status[0] : _GEN_25; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 63:42 71:29]
  assign generateFinalResult_isNaN = _addSub_enable_T_2 ? addSub_status[2] : _GEN_26; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 63:42 72:31]
  assign generateFinalResult_NaNFractionValue = _addSub_enable_T_2 ? addSub_NaNFractionValue : _GEN_27; // @[\\src\\main\\scala\\fpu8\\FPU8Generator.scala 63:42 73:42]
endmodule
